/**************************************************************************/
// Design by Wang Kun Cheng 
// HK416 is my waifu uwu
// Check out the latest version at: https://github.com/I-am-zeroZ/ICLAB_2025_S_pattern
// Feel free to share! The more eyes on this pattern, the more bugs we can squash —
// and the more people get to appreciate how cute HK416 is!
// Welcome to open an issue or even a pull request if you find any bugs or have suggestions.
/**************************************************************************/
`define CYCLE_TIME 20.0
`define PATTERN_NUMBER 10
module PATTERN(
    clk,
    rst_n,
    in_valid,
    in_valid2,
    in_data,
    out_valid,
    out_sad
);
output reg clk, rst_n, in_valid, in_valid2;
output reg [11:0] in_data;
input out_valid;
input out_sad;

//======================================
//      PARAMETERS & VARIABLES
//======================================
integer total_latency;
integer patcount;
integer setcount;
reg [7:0] L0[0:127][0:127];
reg [7:0] L1[0:127][0:127];
reg [7:0] MVinteger_point1[0:63][0:3];  
reg [3:0] MVfraction_point1[0:63][0:3];
reg [7:0] MVinteger_point2[0:63][0:3];  
reg [3:0] MVfraction_point2[0:63][0:3];
reg [15:0] L0_BI_block_result_point1 [0:8][0:7][0:7];
reg [15:0] L1_BI_block_result_point1 [0:8][0:7][0:7];
reg [15:0] L0_BI_block_result_point2 [0:8][0:7][0:7];
reg [15:0] L1_BI_block_result_point2 [0:8][0:7][0:7];
real real_L0_BI_block_result_point1 [0:8][0:7][0:7];
real real_L1_BI_block_result_point1 [0:8][0:7][0:7];
real real_L0_BI_block_result_point2 [0:8][0:7][0:7];
real real_L1_BI_block_result_point2 [0:8][0:7][0:7];
real saved_min_sad_point1, saved_min_sad_point2;
integer saved_search_point_point1, saved_search_point_point2;

reg [55:0] out_sad_got;
reg [55:0] out_sad_golden;


//======================================
//              MAIN
//======================================
initial begin
    total_latency = 0;
    in_valid = 1'b0;
    in_valid2 = 1'b0;
    in_data='x;
    rst_n = 1'b1;
    force clk = 0;
    reset_signal_task;
    for(patcount = 0; patcount < `PATTERN_NUMBER; patcount = patcount + 1) begin
        $display("Pattern %d", patcount);
        generate_testcase; 
        input_task_1;
        @(negedge clk);
        for (setcount = 0; setcount < 64; setcount = setcount + 1) begin
          calculate_ans;
          input_task_2;
          wait_out_valid_task;
          check_ans_task;
        end
    end
    display_pass;
    $finish;
end
//======================================
//              Clock
//======================================
real CYCLE= `CYCLE_TIME;
initial	clk = 0;
always #(CYCLE/2.0) clk = ~clk;

//======================================
//              TASKS
//======================================
task reset_signal_task; 
begin 
  #(0.5);  rst_n=0;
  #(100);  rst_n=1;
  if((out_sad !== 0)||(out_valid !== 0)) 
  begin
    display_fail;
    $display("                    reset_signal_task FAIL                   ");
    $display("**************************************************************");
    $display("*   Output signal should be 0 after initial RESET at %4t     *",$time);
    $display("**************************************************************");
    $finish;
  end
  
  #(3);  release clk;
end 
endtask

integer offset;
integer signed temp;
task generate_testcase;begin
    for(int i=0;i<128;i++)begin
        for(int j=0;j<128;j++)begin
            L0[i][j] = $urandom()%256;
            L1[i][j] = $urandom()%256;
        end
    end
    for (int j=0;j<64;j++) begin
      //MV point1
      for(int i=0;i<4;i++)begin
          MVinteger_point1[j][i] = $urandom()%118; //[0,117]
          MVfraction_point1[j][i] = $urandom()%16; //0~15 (4bit)
      end
      //MV point2
      for(int i=0;i<4;i++)begin
          offset = $urandom()%11-5; //[0,10]-5= [-5,5]
          temp = $signed(MVinteger_point1[j][i]) + offset;
          if(temp < 0)
              temp = 0;
          else if(temp > 117)
              temp = 117;
          MVinteger_point2[j][i] = temp;
          MVfraction_point2[j][i] = $urandom()%16; //0~15 (4bit)  
      end
    end
end
endtask

task input_task_1; 
begin 
    repeat($urandom_range(3,6)-1)@(negedge clk);
    in_valid=1'b1;
    in_valid2=1'b0;
    for(int i=0;i<128;i++)begin
        for(int j=0;j<128;j++)begin
            if(out_valid===1'b1||out_sad!==0)begin
                display_fail;
                $display("\033[0;34mPASS PATTERN NO.%4d,\033[m ",patcount );
                $display("                    input_task FAIL                   ");
                $display("**************************************************************");
                $display("*   The out_valid cannot overlap with in_valid and can rise once for each pattern.  at %4t     *",$time);
                $display("**************************************************************");   
                $finish;
            end
            in_data={L0[i][j],4'bx};
            @(negedge clk);
        end
    end
    for(int i=0;i<128;i++)begin
        for(int j=0;j<128;j++)begin
            if(out_valid===1'b1||out_sad!==0)begin
                display_fail;
                $display("\033[0;34mPASS PATTERN NO.%4d,\033[m ",patcount );
                $display("                    input_task FAIL                   ");
                $display("**************************************************************");
                $display("*   The out_valid cannot overlap with in_valid and can rise once for each pattern.  at %4t     *",$time);
                $display("**************************************************************");   
                $finish;
            end
            in_data={L1[i][j],4'bx};
            @(negedge clk);
        end
    end
    in_valid=1'b0;
    in_data='x;
end
endtask

task input_task_2; 
begin 
    in_valid=1'b0;
    repeat($urandom_range(3,6)-1)@(negedge clk);
    in_valid2=1'b1;
    for(int i=0;i<8;i++)begin
        if(out_valid===1'b1||out_sad!==0)begin
            display_fail;
            $display("\033[0;34mPASS PATTERN NO.%4d,\033[m ",patcount );
            $display("                    input_task FAIL                   ");
            $display("**************************************************************");
            $display("*   The out_valid cannot overlap with in_valid and can rise once for each pattern.  at %4t     *",$time);
            $display("**************************************************************");   
            $finish;
        end
        if(i<4)begin
            in_data={MVinteger_point1[setcount][i],MVfraction_point1[setcount][i]};
        end
        else begin
           in_data={MVinteger_point2[setcount][i-4],MVfraction_point2[setcount][i-4]}; 
        end
        @(negedge clk);
    end

    in_valid2=1'b0;
    in_data='x;
end
endtask

integer wait_val_time;
task wait_out_valid_task;
begin
    wait_val_time = 0;
    while(out_valid!==1'b1) begin
        if(out_sad!==0)begin
            display_fail;
            $display("                   wait_out_valid_task FAIL                   ");
            $display("**************************************************************");
            $display("*    The output signal should be zero when out_valid is low  at %4t     *",$time);
            $display("**************************************************************");           
            $finish;
        end
        wait_val_time=wait_val_time+1;
        if(wait_val_time==1000)begin
            display_fail;
            $display("                    wait_out_valid_task FAIL                   ");
            $display("***************************************************************");
            $display("*         The execution latency are over 1000 cycles.           *");
            $display("***************************************************************");
            repeat(2)@(negedge clk);
            $finish;
        end
        @(negedge clk);
    end
    total_latency = total_latency + wait_val_time;
end
endtask

integer s;
// 搜尋點 offset 陣列 (共 9 個) – L0 用的 offset (dy, dx)
integer L0_dx[0:8], L0_dy[0:8];
// 搜尋點 offset 陣列 (共 9 個) – L1 用的 offset (dy, dx)
integer L1_dx[0:8], L1_dy[0:8];
task calculate_ans; 

  begin
    // 設定 L0 的搜尋點 offset (依照文件中範例)
    L0_dy[0] = 0;  L0_dx[0] = 0;  // Search Pt 0: (0,0)
    L0_dy[1] = 1;  L0_dx[1] = 0;  // Search Pt 1: (1,0)
    L0_dy[2] = 2;  L0_dx[2] = 0;  // Search Pt 2: (2,0)
    L0_dy[3] = 0;  L0_dx[3] = 1;  // Search Pt 3: (0,1)
    L0_dy[4] = 1;  L0_dx[4] = 1;  // Search Pt 4: (1,1)
    L0_dy[5] = 2;  L0_dx[5] = 1;  // Search Pt 5: (2,1)
    L0_dy[6] = 0;  L0_dx[6] = 2;  // Search Pt 6: (0,2)
    L0_dy[7] = 1;  L0_dx[7] = 2;  // Search Pt 7: (1,2)
    L0_dy[8] = 2;  L0_dx[8] = 2;  // Search Pt 8: (2,2)
    
    // 設定 L1 的搜尋點 offset (互補於 L0)
    L1_dy[0] = 2;  L1_dx[0] = 2;  // Search Pt 0: (2,2)
    L1_dy[1] = 1;  L1_dx[1] = 2;  // Search Pt 1: (1,2)
    L1_dy[2] = 0;  L1_dx[2] = 2;  // Search Pt 2: (0,2)
    L1_dy[3] = 2;  L1_dx[3] = 1;  // Search Pt 3: (2,1)
    L1_dy[4] = 1;  L1_dx[4] = 1;  // Search Pt 4: (1,1)
    L1_dy[5] = 0;  L1_dx[5] = 1;  // Search Pt 5: (0,1)
    L1_dy[6] = 2;  L1_dx[6] = 0;  // Search Pt 6: (2,0)
    L1_dy[7] = 1;  L1_dx[7] = 0;  // Search Pt 7: (1,0)
    L1_dy[8] = 0;  L1_dx[8] = 0;  // Search Pt 8: (0,0)
    
    // ====================================================
    // 計算 point1 的 BI 區塊 (共 9 組) 
    // 對於 point1, 
    //   - L0 的 MV 資料: MVinteger_point1[0] 為 MVx, MVinteger_point1[1] 為 MVy
    //   - L1 的 MV 資料: MVinteger_point1[2] 為 MVx, MVinteger_point1[3] 為 MVy
    // ====================================================
    for(s = 0; s < 9; s = s + 1) begin
      // L0 (point1) BI 區塊
      calculate_BI(L0,
                   MVinteger_point1[setcount][0] + L0_dx[s],
                   MVfraction_point1[setcount][0],
                   MVinteger_point1[setcount][1] + L0_dy[s],
                   MVfraction_point1[setcount][1],
                   real_L0_BI_block_result_point1[s]);
                   
      // L1 (point1) BI 區塊
      calculate_BI(L1,
                   MVinteger_point1[setcount][2] + L1_dx[s],
                   MVfraction_point1[setcount][2],
                   MVinteger_point1[setcount][3] + L1_dy[s],
                   MVfraction_point1[setcount][3],
                   real_L1_BI_block_result_point1[s]);
      calculate_sad();
    end
    
    // ====================================================
    // 計算 point2 的 BI 區塊 (共 9 組) 
    // 對於 point2,
    //   - L0 的 MV 資料: MVinteger_point2[0] 為 MVx, MVinteger_point2[1] 為 MVy
    //   - L1 的 MV 資料: MVinteger_point2[2] 為 MVx, MVinteger_point2[3] 為 MVy
    // ====================================================
    for(s = 0; s < 9; s = s + 1) begin
      // L0 (point2) BI 區塊
      calculate_BI(L0,
                   MVinteger_point2[setcount][0] + L0_dx[s],
                   MVfraction_point2[setcount][0],
                   MVinteger_point2[setcount][1] + L0_dy[s],
                   MVfraction_point2[setcount][1],
                   real_L0_BI_block_result_point2[s]);
                   
      // L1 (point2) BI 區塊
      calculate_BI(L1,
                   MVinteger_point2[setcount][2] + L1_dx[s],
                   MVfraction_point2[setcount][2],
                   MVinteger_point2[setcount][3] + L1_dy[s],
                   MVfraction_point2[setcount][3],
                   real_L1_BI_block_result_point2[s]);
      calculate_sad();
    end

  end
endtask


reg [27:0] point1_bits, point2_bits;  
task check_ans_task;
 
begin

  // 連續 56 個 clock 週期擷取序列輸出
  out_sad_got = 56'd0;
  for (int k = 0; k < 56; k = k + 1) begin
    @(posedge clk);
    // 根據 "LSB to MSB" 的描述，先把 out_sad 放在最低 bit，再往高位移
    out_sad_got = {out_sad, out_sad_got[55:1]};
  end

  // 等待 out_valid 拉低 (若 lab 要求)
  while (out_valid === 1'b1) @(negedge clk);

  // 用 function 將 calculate_sad 得到的值 (saved_min_sad_pointX / saved_search_point_pointX)
  // 編碼成 28 bits
  point2_bits = encode_point_and_sad(saved_search_point_point2, saved_min_sad_point2);
  point1_bits = encode_point_and_sad(saved_search_point_point1, saved_min_sad_point1);

  // 圖示中: Output[55:28] => Point2, Output[27:0] => Point1
  // 所以 out_sad_golden = { point2_bits, point1_bits }
  out_sad_golden = {point2_bits, point1_bits};

  // 比對
  if (out_sad_got !== out_sad_golden) begin
    display_fail;
    $display("-----------------------------------------------------");
    $display("  CHECK_ANS FAIL at time %t !!", $time);
    $display("  Got      = %h", out_sad_got);
    $display("  Expected = %h", out_sad_golden);
    $display("-----------------------------------------------------");
    $finish;
  end
  else begin
    // $display("CHECK_ANS PASS at time %t : out_sad = %h", $time, out_sad_got);
  end
end
endtask


task calculate_BI;
  input  [7:0] image [0:127][0:127];
  input  [7:0] MVx_int;    // MV x 整數部分
  input  [3:0] MVx_frac;   // MV x 小數部分 (0~15)
  input  [7:0] MVy_int;    // MV y 整數部分
  input  [3:0] MVy_frac;   // MV y 小數部分 (0~15)
  output real BI_block [0:7][0:7];  // 每個元素為 real 型態
  real x_frac, y_frac;
  real P00, P01, P10, P11;
  real A1, A2, B;
begin
  // 將 4-bit fraction 轉換為 0~1 的比例
  x_frac = MVx_frac / 16.0;
  y_frac = MVy_frac / 16.0;
  
  // 對 8x8 區塊每個點做雙線性插值
  for (int i = 0; i < 8; i = i + 1) begin
    for (int j = 0; j < 8; j = j + 1) begin
      // 取得鄰近的四個像素值，注意影像索引應合法
      P00 = image[MVy_int + i][MVx_int + j];
      P01 = image[MVy_int + i][MVx_int + j + 1];
      P10 = image[MVy_int + i + 1][MVx_int + j];
      P11 = image[MVy_int + i + 1][MVx_int + j + 1];
      
      // 水平插值：先在水平方向算出兩個中間值
      A1 = P00 * (1.0 - x_frac) + P01 * x_frac;
      A2 = P10 * (1.0 - x_frac) + P11 * x_frac;
      
      // 垂直插值：再在垂直方向做插值得到最終值
      B = A1 * (1.0 - y_frac) + A2 * y_frac;
      
      // 將計算結果存入 BI_block 陣列
      BI_block[i][j] = B;
    end
  end
  // calculate_sad(saved_min_sad_point1, saved_search_point_point1,
  //               saved_min_sad_point2, saved_search_point_point2);

end
endtask

// real out_min_sad_point1;
// integer out_min_search_point1;
// real out_min_sad_point2;
// integer out_min_search_point2;
task calculate_sad;
  // output real out_min_sad_point1;
  // output integer out_min_search_point1;
  // output real out_min_sad_point2;
  // output integer out_min_search_point2;
  real sad_point1[0:8];
  real sad_point2[0:8];
  real diff;
  real min_sad1, min_sad2;
  integer min_idx1, min_idx2;
begin
  // 計算 point1 的 SAD 值
  for (int s = 0; s < 9; s = s + 1) begin
    sad_point1[s] = 0.0;
    for (int i = 0; i < 8; i = i + 1) begin
      for (int j = 0; j < 8; j = j + 1) begin
        diff = real_L0_BI_block_result_point1[s][i][j] - real_L1_BI_block_result_point1[s][i][j];
        if (diff < 0)
          diff = -diff;
        sad_point1[s] = sad_point1[s] + diff;
      end
    end
  end
  
  // 計算 point2 的 SAD 值
  for (int s = 0; s < 9; s = s + 1) begin
    sad_point2[s] = 0.0;
    for (int i = 0; i < 8; i = i + 1) begin
      for (int j = 0; j < 8; j = j + 1) begin
        diff = real_L0_BI_block_result_point2[s][i][j] - real_L1_BI_block_result_point2[s][i][j];
        if (diff < 0)
          diff = -diff;
        sad_point2[s] = sad_point2[s] + diff;
      end
    end
  end
  
  // 找出 point1 最小的 SAD 值與搜尋點編號
  min_sad1 = sad_point1[0];
  min_idx1 = 0;
  for (int s = 1; s < 9; s = s + 1) begin
    if (sad_point1[s] < min_sad1) begin
      min_sad1 = sad_point1[s];
      min_idx1 = s;
    end
  end
  
  // 找出 point2 最小的 SAD 值與搜尋點編號
  min_sad2 = sad_point2[0];
  min_idx2 = 0;
  for (int s = 1; s < 9; s = s + 1) begin
    if (sad_point2[s] < min_sad2) begin
      min_sad2 = sad_point2[s];
      min_idx2 = s;
    end
  end
  
  // 將結果以 output 參數輸出，同時更新全域變數
  // out_min_sad_point1 = min_sad1;
  // out_min_search_point1 = min_idx1;
  // out_min_sad_point2 = min_sad2;
  // out_min_search_point2 = min_idx2;
  
  saved_min_sad_point1 = min_sad1;
  saved_search_point_point1 = min_idx1;
  saved_min_sad_point2 = min_sad2;
  saved_search_point_point2 = min_idx2;
  
  // $display("Point1: min SAD = %f at search point %0d", min_sad1, min_idx1);
  // $display("Point2: min SAD = %f at search point %0d", min_sad2, min_idx2);
end
endtask

function [27:0] encode_point_and_sad;
  input integer search_pt;   // 0~8
  input real    sad_value;   // 可能為浮點
  // 若 SAD 可能很大，請檢查 16 bits integer 是否足夠
  reg [15:0] sad_integer;
  reg [7:0]  sad_fraction;
  reg [27:0] out_val;
  real  tmp_real;
begin
  // 1) 取整數部分 (最多支援到 65535)
  //    如果超過範圍要 clamp
  if (sad_value < 0.0)
    sad_value = 0.0;  
  if (sad_value > 65535.0)
    sad_value = 65535.0;
  
  sad_integer = $rtoi(sad_value);  // 截斷或可加 0.5 做四捨五入

  // 2) 取小數部分，轉 8 bits fraction
  //    fraction = (sad_value - sad_integer) * 256
  tmp_real = (sad_value - sad_integer) * 256.0;
  if (tmp_real < 0.0)
    tmp_real = 0.0;
  else if (tmp_real > 255.0)
    tmp_real = 255.0;
  // 四捨五入
  tmp_real = tmp_real + 0.5;  
  sad_fraction = $rtoi(tmp_real);

  // 3) 組合 4 bits search point + 16 bits integer SAD + 8 bits fraction
  out_val = {search_pt[3:0], sad_integer[15:0], sad_fraction[7:0]};
  encode_point_and_sad = out_val;
end
endfunction


task display_fail; begin
    $display("[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m.[0m[38;2;245;245;245m,[0m[38;2;224;224;224m:[0m[38;2;198;198;198m:[0m[38;2;170;170;170m;[0m[38;2;146;146;145m;[0m[38;2;115;115;114m;[0m[38;2;91;91;91m;[0m[38;2;73;73;73m;[0m[38;2;56;56;56m;[0m[38;2;46;46;46m;[0m[38;2;40;40;40m;[0m[38;2;38;38;39mi[0m[38;2;37;37;39mi[0m[38;2;37;37;39mr[0m[38;2;37;37;39mr[0m[38;2;39;38;40mr[0m[38;2;33;33;34mi[0m[38;2;30;30;32mi[0m[38;2;41;41;41mi[0m[38;2;59;59;60mi[0m[38;2;78;79;79mi[0m[38;2;102;102;102m;[0m[38;2;126;126;126m;[0m[38;2;148;148;148m;[0m[38;2;172;172;172m:[0m[38;2;195;195;194m:[0m[38;2;214;214;214m:[0m[38;2;232;232;232m,[0m[38;2;245;245;245m,[0m[38;2;255;255;255m.[0m[38;2;255;255;255m.[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m");
    $display("[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;247;247;246m.[0m[38;2;207;207;207m:[0m[38;2;153;153;153m;[0m[38;2;95;95;95m;[0m[38;2;55;55;56m;[0m[38;2;37;37;38m;[0m[38;2;28;28;30mi[0m[38;2;27;27;29mr[0m[38;2;29;30;33mr[0m[38;2;36;36;40ms[0m[38;2;42;42;47mX[0m[38;2;49;50;55mA[0m[38;2;57;57;62m2[0m[38;2;61;61;67m2[0m[38;2;67;67;74m5[0m[38;2;72;72;79m3[0m[38;2;75;75;83m3[0m[38;2;78;78;86m3[0m[38;2;79;79;87m3[0m[38;2;80;80;87m3[0m[38;2;79;79;87m3[0m[38;2;75;75;83m3[0m[38;2;71;71;78m5[0m[38;2;68;68;75m5[0m[38;2;63;64;70m5[0m[38;2;56;57;62m2[0m[38;2;52;52;57m2[0m[38;2;46;47;51mA[0m[38;2;41;42;46mX[0m[38;2;38;38;41ms[0m[38;2;38;38;40mi[0m[38;2;40;40;41m;[0m[38;2;49;49;50m:[0m[38;2;70;70;69m:[0m[38;2;107;107;107m;[0m[38;2;151;151;151m;[0m[38;2;209;209;209m:[0m[38;2;251;251;251m,[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m");
    $display("[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;242;242;242m,[0m[38;2;202;202;203m;[0m[38;2;149;149;151ms[0m[38;2;90;90;93mA[0m[38;2;60;60;65m2[0m[38;2;52;53;58m2[0m[38;2;57;57;64m2[0m[38;2;65;65;71m5[0m[38;2;73;73;81m3[0m[38;2;79;79;86m3[0m[38;2;82;82;90mh[0m[38;2;84;84;92mh[0m[38;2;85;85;93mh[0m[38;2;85;85;93mh[0m[38;2;85;85;93mh[0m[38;2;84;84;93mh[0m[38;2;84;84;92mh[0m[38;2;83;83;92mh[0m[38;2;83;83;91mh[0m[38;2;83;83;91mh[0m[38;2;82;82;91mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;83;83;91mh[0m[38;2;83;83;91mh[0m[38;2;83;83;91mh[0m[38;2;84;84;92mh[0m[38;2;84;84;92mh[0m[38;2;84;84;93mh[0m[38;2;84;84;93mh[0m[38;2;84;84;92mh[0m[38;2;82;82;91mh[0m[38;2;78;78;86m3[0m[38;2;70;69;77m5[0m[38;2;56;56;62m2[0m[38;2;39;39;44mX[0m[38;2;20;20;24mi[0m[38;2;7;8;9m:[0m[38;2;14;14;15m:[0m[38;2;66;66;66m;[0m[38;2;154;154;154mi[0m[38;2;227;227;227m:[0m[38;2;255;255;255m.[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m");
    $display("[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m.[0m[38;2;241;241;241m,[0m[38;2;189;189;189m;[0m[38;2;134;134;136mX[0m[38;2;95;95;99m5[0m[38;2;75;76;82m3[0m[38;2;73;73;82mh[0m[38;2;78;78;86mh[0m[38;2;83;83;91mh[0m[38;2;84;84;92mh[0m[38;2;84;84;92mh[0m[38;2;83;83;92mh[0m[38;2;83;83;91mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;91mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;91mh[0m[38;2;83;83;91mh[0m[38;2;84;84;92mh[0m[38;2;85;85;93mh[0m[38;2;83;84;92mh[0m[38;2;78;78;86m3[0m[38;2;62;63;70m2[0m[38;2;33;33;36ms[0m[38;2;10;11;12m;[0m[38;2;29;29;29m:[0m[38;2;97;97;97m;[0m[38;2;183;183;182m;[0m[38;2;247;247;247m,[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m");
    $display("[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;249;249;249m,[0m[38;2;196;196;196m:[0m[38;2;124;125;125mi[0m[38;2;77;78;81mX[0m[38;2;63;63;69m5[0m[38;2;67;67;75m3[0m[38;2;72;72;80m3[0m[38;2;76;76;84m3[0m[38;2;82;83;91mh[0m[38;2;83;83;91mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;81;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;84;84;92mh[0m[38;2;85;85;93mh[0m[38;2;85;85;93mh[0m[38;2;83;83;91mh[0m[38;2;82;82;90mh[0m[38;2;81;81;89mh[0m[38;2;81;81;89mh[0m[38;2;81;81;89mh[0m[38;2;82;82;90mh[0m[38;2;83;83;91mh[0m[38;2;84;84;92mh[0m[38;2;85;85;93mh[0m[38;2;84;84;93mh[0m[38;2;84;84;92mh[0m[38;2;83;83;91mh[0m[38;2;83;82;91mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;83;83;91mh[0m[38;2;84;84;92mh[0m[38;2;85;85;93mh[0m[38;2;77;77;85m3[0m[38;2;53;54;60mA[0m[38;2;21;22;25mi[0m[38;2;8;8;9m:[0m[38;2;55;55;55m;[0m[38;2;154;154;154mi[0m[38;2;237;237;237m:[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;252;252;252m,[0m[38;2;220;220;219m:[0m[38;2;190;190;190m:[0m[38;2;185;185;185m:[0m[38;2;208;208;208m:[0m[38;2;243;243;243m,[0m[38;2;255;255;255m.[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m");
    $display("[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m.[0m[38;2;225;225;225m:[0m[38;2;151;151;151m;[0m[38;2;63;63;63m;[0m[38;2;8;8;8m,[0m[38;2;9;9;11m;[0m[38;2;19;19;22m;[0m[38;2;19;19;21m;[0m[38;2;15;15;17m:[0m[38;2;10;10;12m,[0m[38;2;12;12;13m:[0m[38;2;29;30;33mi[0m[38;2;71;72;79m5[0m[38;2;84;84;92mh[0m[38;2;83;83;91mh[0m[38;2;83;83;91mh[0m[38;2;83;82;91mh[0m[38;2;83;83;91mh[0m[38;2;82;82;90mh[0m[38;2;65;65;71m5[0m[38;2;45;45;49mX[0m[38;2;33;34;36mr[0m[38;2;21;22;24m;[0m[38;2;16;17;19m:[0m[38;2;14;14;16m:[0m[38;2;14;13;14m:[0m[38;2;14;15;17m:[0m[38;2;16;16;18m:[0m[38;2;19;19;22m;[0m[38;2;32;31;35mr[0m[38;2;46;47;51mX[0m[38;2;57;58;63m2[0m[38;2;68;68;74m5[0m[38;2;76;76;83m3[0m[38;2;81;81;89mh[0m[38;2;83;83;92mh[0m[38;2;85;85;93mh[0m[38;2;85;85;93mh[0m[38;2;84;84;93mh[0m[38;2;84;84;92mh[0m[38;2;83;83;91mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;83;83;91mh[0m[38;2;84;85;93mh[0m[38;2;83;83;91mh[0m[38;2;67;67;74m5[0m[38;2;30;30;33mr[0m[38;2;5;4;5m:[0m[38;2;48;48;47m;[0m[38;2;153;153;153mi[0m[38;2;242;242;242m:[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;247;247;247m,[0m[38;2;164;164;163mi[0m[38;2;66;66;66m;[0m[38;2;28;28;29m;[0m[38;2;43;44;46mX[0m[38;2;49;50;52mA[0m[38;2;33;33;34mr[0m[38;2;45;44;45m:[0m[38;2;114;114;114m;[0m[38;2;207;207;207m;[0m[38;2;255;255;255m.[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m");
    $display("[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m,[0m[38;2;222;222;222m:[0m[38;2;160;160;160m;[0m[38;2;85;85;84m:[0m[38;2;24;24;24m:[0m[38;2;5;5;6m:[0m[38;2;24;24;26mi[0m[38;2;54;54;57mA[0m[38;2;81;81;86m3[0m[38;2;68;68;73m5[0m[38;2;53;54;59mA[0m[38;2;49;49;53mX[0m[38;2;8;8;8m,[0m[38;2;13;13;13m:[0m[38;2;2;2;2m.[0m[38;2;32;32;35mr[0m[38;2;74;74;81m3[0m[38;2;76;76;83m3[0m[38;2;78;78;86m3[0m[38;2;80;81;89mh[0m[38;2;76;77;85m3[0m[38;2;33;34;38mr[0m[38;2;3;3;3m.[0m[38;2;0;0;0m [0m[38;2;0;0;0m [0m[38;2;66;66;70m5[0m[38;2;88;87;93mh[0m[38;2;77;76;81m3[0m[38;2;64;64;70m2[0m[38;2;51;51;54mA[0m[38;2;38;37;39ms[0m[38;2;28;28;30mi[0m[38;2;15;15;16m:[0m[38;2;8;8;8m,[0m[38;2;2;2;2m.[0m[38;2;1;1;1m.[0m[38;2;4;5;6m.[0m[38;2;12;12;13m:[0m[38;2;22;23;25m;[0m[38;2;34;34;37mr[0m[38;2;47;47;51mX[0m[38;2;59;59;65m2[0m[38;2;70;70;77m5[0m[38;2;77;77;85m3[0m[38;2;82;82;90mh[0m[38;2;84;84;93mh[0m[38;2;85;85;93mh[0m[38;2;84;84;92mh[0m[38;2;83;83;91mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;83;83;91mh[0m[38;2;82;82;90mh[0m[38;2;66;65;72m5[0m[38;2;26;26;29mi[0m[38;2;3;3;3m,[0m[38;2;54;54;54m;[0m[38;2;172;172;172mi[0m[38;2;252;252;252m,[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m.[0m[38;2;205;205;205m;[0m[38;2;70;70;69m;[0m[38;2;10;10;11m:[0m[38;2;84;85;89mM[0m[38;2;180;182;188m&[0m[38;2;224;227;233m@[0m[38;2;229;232;237m@[0m[38;2;205;207;212m@[0m[38;2;139;141;145m#[0m[38;2;49;49;51mA[0m[38;2;16;16;16m:[0m[38;2;105;105;105m;[0m[38;2;222;222;222m;[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m");
    $display("[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m.[0m[38;2;222;222;222m:[0m[38;2;145;145;145mi[0m[38;2;68;68;68m:[0m[38;2;20;20;20m:[0m[38;2;22;22;24mr[0m[38;2;67;67;73m3[0m[38;2;115;115;125mG[0m[38;2;144;142;153m9[0m[38;2;162;161;174mB[0m[38;2;171;170;184mB[0m[38;2;175;174;189m&[0m[38;2;122;122;131mS[0m[38;2;78;79;87m3[0m[38;2;66;66;71m5[0m[38;2;11;11;11m,[0m[38;2;12;12;12m,[0m[38;2;9;9;9m,[0m[38;2;3;4;4m.[0m[38;2;14;14;16m:[0m[38;2;16;16;17m:[0m[38;2;16;16;18m:[0m[38;2;18;18;21m;[0m[38;2;14;15;17m:[0m[38;2;0;0;0m [0m[38;2;0;0;0m [0m[38;2;0;0;0m [0m[38;2;47;47;49mX[0m[38;2;163;162;175mB[0m[38;2;177;176;190m&[0m[38;2;175;174;188m&[0m[38;2;174;173;187mB[0m[38;2;171;170;184mB[0m[38;2;168;167;180mB[0m[38;2;164;163;176mB[0m[38;2;154;153;165m9[0m[38;2;147;146;157m9[0m[38;2;132;130;141m#[0m[38;2;115;114;122mG[0m[38;2;92;92;98mM[0m[38;2;69;69;74m5[0m[38;2;46;45;48mX[0m[38;2;24;24;26mi[0m[38;2;8;8;8m,[0m[38;2;0;0;0m [0m[38;2;0;0;0m [0m[38;2;8;8;9m,[0m[38;2;19;20;22m;[0m[38;2;34;34;37mr[0m[38;2;50;50;55mA[0m[38;2;65;65;72m5[0m[38;2;77;78;85m3[0m[38;2;83;83;91mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;80;80;88m3[0m[38;2;78;78;86m3[0m[38;2;80;80;87m3[0m[38;2;83;83;91mh[0m[38;2;89;89;97mh[0m[38;2;99;98;106mM[0m[38;2;111;111;120mG[0m[38;2;120;121;130mS[0m[38;2;75;75;81m3[0m[38;2;19;18;21m;[0m[38;2;4;4;4m,[0m[38;2;93;93;93mi[0m[38;2;224;224;224m;[0m[38;2;255;255;255m [0m[38;2;254;254;254m,[0m[38;2;159;159;159mr[0m[38;2;20;20;20m:[0m[38;2;33;34;36ms[0m[38;2;167;168;173mB[0m[38;2;238;241;246m@[0m[38;2;241;245;249m@[0m[38;2;237;240;245m@[0m[38;2;237;240;245m@[0m[38;2;239;242;247m@[0m[38;2;243;247;252m@[0m[38;2;228;230;235m@[0m[38;2;140;140;144m#[0m[38;2;20;20;21mi[0m[38;2;34;34;34m:[0m[38;2;176;176;176mr[0m[38;2;255;255;255m.[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m");
    $display("[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;227;227;227m:[0m[38;2;113;113;113mi[0m[38;2;23;23;23m:[0m[38;2;7;7;8m:[0m[38;2;58;57;61m2[0m[38;2;116;116;124mG[0m[38;2;158;158;170mB[0m[38;2;174;173;187mB[0m[38;2;175;173;188m&[0m[38;2;173;172;186mB[0m[38;2;172;171;185mB[0m[38;2;172;171;185mB[0m[38;2;173;173;188mB[0m[38;2;123;123;133mS[0m[38;2;77;78;86m3[0m[38;2;69;71;78m5[0m[38;2;15;15;17m:[0m[38;2;11;11;10m,[0m[38;2;10;9;9m,[0m[38;2;15;16;18m:[0m[38;2;60;61;67m2[0m[38;2;64;65;71m2[0m[38;2;62;63;69m2[0m[38;2;45;46;51mX[0m[38;2;3;3;4m.[0m[38;2;0;0;0m [0m[38;2;0;0;0m [0m[38;2;10;10;11m,[0m[38;2;125;124;133mS[0m[38;2;173;172;186mB[0m[38;2;169;168;182mB[0m[38;2;169;168;182mB[0m[38;2;169;168;182mB[0m[38;2;169;168;183mB[0m[38;2;170;169;183mB[0m[38;2;170;169;183mB[0m[38;2;171;170;185mB[0m[38;2;172;171;185mB[0m[38;2;173;172;187mB[0m[38;2;174;173;188m&[0m[38;2;175;174;189m&[0m[38;2;174;173;187mB[0m[38;2;170;169;182mB[0m[38;2;161;160;173mB[0m[38;2;144;144;155m9[0m[38;2;120;120;129mS[0m[38;2;87;87;93mh[0m[38;2;40;40;42ms[0m[38;2;9;9;9m,[0m[38;2;0;0;0m [0m[38;2;0;0;0m [0m[38;2;2;2;2m.[0m[38;2;13;13;14m:[0m[38;2;43;44;47mX[0m[38;2;81;81;89mh[0m[38;2;82;81;89mh[0m[38;2;102;102;109mH[0m[38;2;136;136;148m#[0m[38;2;150;151;164m9[0m[38;2;162;163;176mB[0m[38;2;172;173;188mB[0m[38;2;181;181;197m&[0m[38;2;186;186;203m&[0m[38;2;189;190;207m&[0m[38;2;156;156;168m9[0m[38;2;85;85;91mh[0m[38;2;44;45;49mX[0m[38;2;1;1;1m,[0m[38;2;49;49;49mi[0m[38;2;179;179;179mr[0m[38;2;120;120;120mr[0m[38;2;5;5;6m,[0m[38;2;64;64;67m5[0m[38;2;202;204;210m@[0m[38;2;242;245;250m@[0m[38;2;236;239;244m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;237;240;245m@[0m[38;2;243;246;251m@[0m[38;2;190;192;197m&[0m[38;2;50;50;53mA[0m[38;2;10;10;9m,[0m[38;2;136;136;136mr[0m[38;2;247;247;247m,[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m");
    $display("[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;245;245;245m,[0m[38;2;150;150;150mi[0m[38;2;40;40;40m;[0m[38;2;1;1;2m,[0m[38;2;77;77;83m3[0m[38;2;145;144;155m9[0m[38;2;173;172;186mB[0m[38;2;176;175;189m&[0m[38;2;174;173;187mB[0m[38;2;175;173;188m&[0m[38;2;175;174;188m&[0m[38;2;172;171;185mB[0m[38;2;164;163;177mB[0m[38;2;152;152;164m9[0m[38;2;134;134;144m#[0m[38;2;90;90;96mM[0m[38;2;65;66;72m5[0m[38;2;57;58;64m2[0m[38;2;12;12;14m:[0m[38;2;8;8;7m,[0m[38;2;8;8;8m,[0m[38;2;6;6;6m,[0m[38;2;18;18;20m;[0m[38;2;22;22;24m;[0m[38;2;27;27;30mi[0m[38;2;20;20;22m;[0m[38;2;0;0;0m [0m[38;2;0;0;0m [0m[38;2;0;0;0m [0m[38;2;65;65;69m2[0m[38;2;173;172;186mB[0m[38;2;174;172;187mB[0m[38;2;170;169;183mB[0m[38;2;169;168;182mB[0m[38;2;169;168;182mB[0m[38;2;169;168;182mB[0m[38;2;169;168;182mB[0m[38;2;169;168;182mB[0m[38;2;169;168;182mB[0m[38;2;169;168;182mB[0m[38;2;169;168;182mB[0m[38;2;169;168;182mB[0m[38;2;169;168;182mB[0m[38;2;169;168;182mB[0m[38;2;170;169;183mB[0m[38;2;171;170;184mB[0m[38;2;172;171;186mB[0m[38;2;174;173;188m&[0m[38;2;176;175;188m&[0m[38;2;124;123;131mS[0m[38;2;71;72;79m5[0m[38;2;63;64;71m2[0m[38;2;42;42;46ms[0m[38;2;4;4;4m.[0m[38;2;0;0;0m [0m[38;2;5;5;5m.[0m[38;2;55;56;62mA[0m[38;2;81;81;89mh[0m[38;2;100;100;107mH[0m[38;2;168;169;182mB[0m[38;2;191;192;209m&[0m[38;2;188;188;205m&[0m[38;2;187;187;204m&[0m[38;2;186;187;204m&[0m[38;2;186;186;203m&[0m[38;2;186;186;203m&[0m[38;2;187;187;204m&[0m[38;2;138;139;151m#[0m[38;2;86;86;93mh[0m[38;2;58;58;64m2[0m[38;2;7;7;8m,[0m[38;2;3;3;3m,[0m[38;2;2;2;3m,[0m[38;2;98;99;102mM[0m[38;2;222;225;230m@[0m[38;2;240;243;248m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;241;244;249m@[0m[38;2;215;217;222m@[0m[38;2;78;79;83m3[0m[38;2;0;0;1m,[0m[38;2;102;102;101mr[0m[38;2;240;240;240m:[0m[38;2;255;255;255m [0m");
    $display("[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;251;251;251m,[0m[38;2;130;130;130ms[0m[38;2;2;2;2m:[0m[38;2;1;1;2m.[0m[38;2;92;91;98mM[0m[38;2;177;176;190m&[0m[38;2;179;178;192m&[0m[38;2;172;171;185mB[0m[38;2;162;161;174mB[0m[38;2;144;143;155m9[0m[38;2;116;116;125mG[0m[38;2;85;85;92mh[0m[38;2;57;57;61mA[0m[38;2;34;34;37mr[0m[38;2;18;18;20m;[0m[38;2;8;8;8m,[0m[38;2;5;5;5m.[0m[38;2;7;8;8m,[0m[38;2;7;7;8m,[0m[38;2;9;9;10m,[0m[38;2;15;15;19m:[0m[38;2;24;25;30mi[0m[38;2;25;26;32mi[0m[38;2;22;24;29mi[0m[38;2;20;22;27m;[0m[38;2;18;19;24m;[0m[38;2;13;14;18m:[0m[38;2;8;9;10m,[0m[38;2;1;1;1m.[0m[38;2;0;0;0m [0m[38;2;47;47;50mX[0m[38;2;107;107;115mH[0m[38;2;143;142;154m9[0m[38;2;166;165;179mB[0m[38;2;174;173;188m&[0m[38;2;175;174;188m&[0m[38;2;172;171;185mB[0m[38;2;170;169;183mB[0m[38;2;169;168;182mB[0m[38;2;169;168;182mB[0m[38;2;169;168;182mB[0m[38;2;169;168;182mB[0m[38;2;169;168;182mB[0m[38;2;169;168;182mB[0m[38;2;169;168;182mB[0m[38;2;169;168;182mB[0m[38;2;169;168;182mB[0m[38;2;169;168;182mB[0m[38;2;169;168;182mB[0m[38;2;170;169;182mB[0m[38;2;123;123;130mS[0m[38;2;76;77;85m3[0m[38;2;79;80;88m3[0m[38;2;69;69;76m5[0m[38;2;11;10;11m,[0m[38;2;0;0;0m [0m[38;2;0;0;0m [0m[38;2;26;27;32mi[0m[38;2;73;74;81m3[0m[38;2;80;80;88m3[0m[38;2;103;102;109mH[0m[38;2;172;173;187mB[0m[38;2;187;188;205m&[0m[38;2;185;186;202m&[0m[38;2;185;186;203m&[0m[38;2;186;186;203m&[0m[38;2;186;187;204m&[0m[38;2;188;188;206m&[0m[38;2;188;189;206m&[0m[38;2;141;143;155m9[0m[38;2;112;112;121mG[0m[38;2;118;118;127mG[0m[38;2;39;39;41ms[0m[38;2;1;2;2m.[0m[38;2;128;130;135mS[0m[38;2;239;242;247m@[0m[38;2;236;239;244m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;240;243;248m@[0m[38;2;224;227;232m@[0m[38;2;93;94;97mM[0m[38;2;0;0;0m.[0m[38;2;95;95;96mr[0m[38;2;240;240;240m:[0m");
    $display("[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;241;241;241m:[0m[38;2;67;67;67ms[0m[38;2;0;0;0m [0m[38;2;30;30;31mi[0m[38;2;126;126;135mS[0m[38;2;113;112;121mG[0m[38;2;80;79;85m3[0m[38;2;51;51;55mA[0m[38;2;26;26;28mi[0m[38;2;6;6;7m,[0m[38;2;0;0;0m [0m[38;2;0;0;0m [0m[38;2;0;0;0m [0m[38;2;0;0;0m [0m[38;2;2;2;2m.[0m[38;2;3;4;4m.[0m[38;2;4;4;5m.[0m[38;2;7;7;7m,[0m[38;2;9;9;10m,[0m[38;2;12;12;14m:[0m[38;2;13;14;16m:[0m[38;2;14;15;18m:[0m[38;2;17;18;22m;[0m[38;2;19;20;24m;[0m[38;2;21;22;28m;[0m[38;2;22;24;30mi[0m[38;2;24;26;32mi[0m[38;2;24;26;33mi[0m[38;2;19;20;25m;[0m[38;2;10;11;13m,[0m[38;2;2;2;3m.[0m[38;2;0;0;0m [0m[38;2;9;9;9m,[0m[38;2;36;36;38mr[0m[38;2;73;73;78m5[0m[38;2;114;113;122mG[0m[38;2;148;146;158m9[0m[38;2;167;166;180mB[0m[38;2;174;173;188m&[0m[38;2;174;173;188m&[0m[38;2;172;171;186mB[0m[38;2;171;170;184mB[0m[38;2;170;169;183mB[0m[38;2;169;168;182mB[0m[38;2;169;168;182mB[0m[38;2;169;168;182mB[0m[38;2;169;168;182mB[0m[38;2;169;168;182mB[0m[38;2;169;168;182mB[0m[38;2;170;169;182mB[0m[38;2;119;120;126mG[0m[38;2;74;75;83m3[0m[38;2;77;78;86m3[0m[38;2;65;66;73m5[0m[38;2;9;9;10m,[0m[38;2;0;0;0m [0m[38;2;0;0;1m.[0m[38;2;23;24;29mi[0m[38;2;64;65;71m2[0m[38;2;81;81;88mh[0m[38;2;77;76;84m3[0m[38;2;117;117;125mG[0m[38;2;178;179;195m&[0m[38;2;187;188;205m&[0m[38;2;188;189;206m&[0m[38;2;186;187;203m&[0m[38;2;180;180;196m&[0m[38;2;169;169;183mB[0m[38;2;161;162;175mB[0m[38;2;182;182;198m&[0m[38;2;187;188;204m&[0m[38;2;191;192;210m&[0m[38;2;157;158;169mB[0m[38;2;41;41;43ms[0m[38;2;8;8;9m,[0m[38;2;146;147;152m9[0m[38;2;238;241;246m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;239;242;247m@[0m[38;2;225;227;233m@[0m[38;2;94;94;97mM[0m[38;2;0;0;0m.[0m[38;2;102;102;102mr[0m");
    $display("[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;237;237;237m;[0m[38;2;55;55;55mr[0m[38;2;0;0;0m [0m[38;2;6;6;6m,[0m[38;2;5;6;6m.[0m[38;2;0;0;0m [0m[38;2;4;4;4m.[0m[38;2;13;13;15m:[0m[38;2;25;25;29mi[0m[38;2;36;36;40mr[0m[38;2;46;46;50mX[0m[38;2;52;52;57mA[0m[38;2;56;56;61mA[0m[38;2;59;59;65m2[0m[38;2;62;62;69m2[0m[38;2;64;64;70m2[0m[38;2;65;65;71m5[0m[38;2;66;65;71m5[0m[38;2;66;66;72m5[0m[38;2;66;66;72m5[0m[38;2;65;65;71m5[0m[38;2;64;64;69m2[0m[38;2;63;63;69m2[0m[38;2;63;63;69m2[0m[38;2;60;60;66m2[0m[38;2;57;58;63m2[0m[38;2;54;53;58mA[0m[38;2;42;42;47ms[0m[38;2;30;30;34mr[0m[38;2;23;23;26m;[0m[38;2;16;17;19m:[0m[38;2;12;13;16m:[0m[38;2;9;9;12m,[0m[38;2;3;4;5m.[0m[38;2;0;0;0m [0m[38;2;0;0;0m [0m[38;2;12;12;12m:[0m[38;2;40;40;43ms[0m[38;2;77;77;84m3[0m[38;2;113;114;123mG[0m[38;2;141;141;152m#[0m[38;2;160;159;172mB[0m[38;2;168;167;181mB[0m[38;2;172;171;185mB[0m[38;2;172;171;186mB[0m[38;2;172;171;185mB[0m[38;2;171;170;184mB[0m[38;2;170;169;183mB[0m[38;2;169;168;182mB[0m[38;2;168;168;182mB[0m[38;2;113;114;121mG[0m[38;2;74;75;83m3[0m[38;2;77;78;87m3[0m[38;2;65;66;73m5[0m[38;2;9;9;10m,[0m[38;2;0;0;0m [0m[38;2;4;4;5m.[0m[38;2;29;30;36mr[0m[38;2;71;71;78m5[0m[38;2;103;103;111mH[0m[38;2;120;119;129mS[0m[38;2;148;148;159m9[0m[38;2;181;181;197m&[0m[38;2;172;173;188mB[0m[38;2;129;129;139mS[0m[38;2;111;111;120mG[0m[38;2;98;98;106mM[0m[38;2;87;87;94mh[0m[38;2;82;81;89mh[0m[38;2;128;128;138mS[0m[38;2;185;186;202m&[0m[38;2;186;186;203m&[0m[38;2;190;190;208m&[0m[38;2;159;159;173mB[0m[38;2;40;40;43ms[0m[38;2;23;23;24m;[0m[38;2;186;188;194m&[0m[38;2;239;242;247m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;239;242;247m@[0m[38;2;222;225;230m@[0m[38;2;78;78;81m3[0m[38;2;1;1;1m.[0m");
    $display("[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m.[0m[38;2;237;237;237m,[0m[38;2;197;197;197m:[0m[38;2;145;145;145m;[0m[38;2;87;87;87mi[0m[38;2;15;15;16m:[0m[38;2;21;21;24m;[0m[38;2;42;42;46ms[0m[38;2;59;59;65m2[0m[38;2;70;71;77m5[0m[38;2;78;78;86m3[0m[38;2;84;84;92mh[0m[38;2;86;86;95mh[0m[38;2;87;87;95mh[0m[38;2;87;87;95mh[0m[38;2;86;86;95mh[0m[38;2;86;86;94mh[0m[38;2;85;85;93mh[0m[38;2;84;84;93mh[0m[38;2;84;84;92mh[0m[38;2;84;84;92mh[0m[38;2;84;84;92mh[0m[38;2;84;84;92mh[0m[38;2;84;84;92mh[0m[38;2;84;84;92mh[0m[38;2;84;84;92mh[0m[38;2;84;84;92mh[0m[38;2;84;84;92mh[0m[38;2;84;84;92mh[0m[38;2;84;84;93mh[0m[38;2;85;85;93mh[0m[38;2;84;84;92mh[0m[38;2;82;81;89mh[0m[38;2;76;75;82m3[0m[38;2;65;65;71m5[0m[38;2;51;51;56mA[0m[38;2;34;34;38mr[0m[38;2;19;19;21m;[0m[38;2;9;9;11m,[0m[38;2;3;4;4m.[0m[38;2;0;0;0m [0m[38;2;0;0;0m [0m[38;2;0;0;0m [0m[38;2;0;0;0m [0m[38;2;13;13;14m:[0m[38;2;39;40;43ms[0m[38;2;72;73;78m5[0m[38;2;105;105;112mH[0m[38;2;129;129;139mS[0m[38;2;146;145;156m9[0m[38;2;157;156;168m9[0m[38;2;165;164;177mB[0m[38;2;171;169;183mB[0m[38;2;170;170;184mB[0m[38;2;105;106;117mH[0m[38;2;74;75;82m3[0m[38;2;77;78;87m3[0m[38;2;64;66;73m5[0m[38;2;8;9;10m,[0m[38;2;0;0;0m [0m[38;2;43;43;47ms[0m[38;2;151;151;163m9[0m[38;2;172;172;187mB[0m[38;2;183;183;199m&[0m[38;2;188;188;205m&[0m[38;2;188;189;206m&[0m[38;2;188;188;205m&[0m[38;2;168;169;183mB[0m[38;2;93;93;100mM[0m[38;2;77;77;85m3[0m[38;2;81;81;89mh[0m[38;2;83;83;91mh[0m[38;2;82;82;90mh[0m[38;2;87;86;93mh[0m[38;2;158;158;170mB[0m[38;2;193;194;211m&[0m[38;2;189;190;207m&[0m[38;2;169;169;184mB[0m[38;2;81;82;88mh[0m[38;2;0;0;0m [0m[38;2;88;89;92mh[0m[38;2;232;234;240m@[0m[38;2;236;239;244m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;240;243;248m@[0m[38;2;202;205;210m@[0m[38;2;50;50;52mX[0m");
    $display("[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m.[0m[38;2;242;242;242m,[0m[38;2;195;195;195m;[0m[38;2;134;134;134m;[0m[38;2;77;77;77m;[0m[38;2;33;33;33m:[0m[38;2;8;8;8m:[0m[38;2;2;2;4m:[0m[38;2;12;12;15m;[0m[38;2;34;34;37mr[0m[38;2;45;45;48mX[0m[38;2;45;45;49mX[0m[38;2;45;45;48mX[0m[38;2;45;44;48mX[0m[38;2;46;45;49mX[0m[38;2;49;49;54mX[0m[38;2;54;55;60mA[0m[38;2;58;58;63m2[0m[38;2;63;63;69m2[0m[38;2;69;70;76m5[0m[38;2;75;75;82m3[0m[38;2;79;80;87m3[0m[38;2;83;83;91mh[0m[38;2;85;85;93mh[0m[38;2;85;85;93mh[0m[38;2;84;84;92mh[0m[38;2;83;83;91mh[0m[38;2;83;83;91mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;83;83;91mh[0m[38;2;84;84;92mh[0m[38;2;85;85;93mh[0m[38;2;83;84;91mh[0m[38;2;78;78;85m3[0m[38;2;65;66;72m5[0m[38;2;50;50;55mA[0m[38;2;35;35;38mr[0m[38;2;20;20;22m;[0m[38;2;8;8;9m,[0m[38;2;2;2;2m.[0m[38;2;0;0;0m [0m[38;2;0;0;0m [0m[38;2;0;0;0m [0m[38;2;7;8;8m,[0m[38;2;27;27;29mi[0m[38;2;50;50;55mA[0m[38;2;72;73;80m3[0m[38;2;92;92;99mM[0m[38;2;108;108;117mH[0m[38;2;121;121;131mS[0m[38;2;91;92;100mM[0m[38;2;75;76;84m3[0m[38;2;78;79;87m3[0m[38;2;54;55;61mA[0m[38;2;3;4;4m.[0m[38;2;0;0;0m [0m[38;2;40;40;45ms[0m[38;2;165;166;180mB[0m[38;2;191;192;209m&[0m[38;2;186;186;203m&[0m[38;2;185;186;203m&[0m[38;2;185;186;202m&[0m[38;2;185;186;203m&[0m[38;2;188;188;205m&[0m[38;2;140;142;154m#[0m[38;2;79;79;87m3[0m[38;2;72;72;80m5[0m[38;2;64;65;72m5[0m[38;2;55;55;62mA[0m[38;2;41;43;50mX[0m[38;2;80;81;89mh[0m[38;2;128;128;139mS[0m[38;2;65;65;71m5[0m[38;2;25;25;27mi[0m[38;2;17;18;19m:[0m[38;2;1;1;1m.[0m[38;2;34;34;36mr[0m[38;2;200;202;208m@[0m[38;2;239;242;247m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;238;241;246m@[0m[38;2;178;179;185m&[0m");
    $display("[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;241;241;241m:[0m[38;2;185;185;185m;[0m[38;2;107;107;107mi[0m[38;2;42;42;42m:[0m[38;2;3;3;3m,[0m[38;2;0;0;0m.[0m[38;2;0;0;0m [0m[38;2;0;0;0m.[0m[38;2;8;8;9m,[0m[38;2;11;11;11m,[0m[38;2;18;20;23m;[0m[38;2;48;53;61mA[0m[38;2;51;57;65mA[0m[38;2;52;57;66mA[0m[38;2;52;58;66mA[0m[38;2;51;56;65mA[0m[38;2;52;57;66mA[0m[38;2;34;38;43ms[0m[38;2;23;25;30mi[0m[38;2;32;35;41mr[0m[38;2;24;26;31mi[0m[38;2;19;21;23m;[0m[38;2;17;17;19m:[0m[38;2;18;18;20m;[0m[38;2;23;23;24m;[0m[38;2;33;32;35mr[0m[38;2;46;46;50mX[0m[38;2;60;59;65m2[0m[38;2;70;71;77m5[0m[38;2;79;79;87m3[0m[38;2;84;84;92mh[0m[38;2;85;85;93mh[0m[38;2;84;84;92mh[0m[38;2;83;83;91mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;83;83;91mh[0m[38;2;84;84;92mh[0m[38;2;85;85;93mh[0m[38;2;84;84;93mh[0m[38;2;81;81;89mh[0m[38;2;72;72;79m5[0m[38;2;59;59;65m2[0m[38;2;42;43;47ms[0m[38;2;23;23;25m;[0m[38;2;6;7;7m,[0m[38;2;0;0;0m [0m[38;2;0;0;0m [0m[38;2;0;0;0m [0m[38;2;6;6;7m,[0m[38;2;21;21;23m;[0m[38;2;42;42;46ms[0m[38;2;62;62;69m2[0m[38;2;76;76;84m3[0m[38;2;77;78;86m3[0m[38;2;79;80;88m3[0m[38;2;39;40;44ms[0m[38;2;0;0;0m [0m[38;2;2;2;3m.[0m[38;2;22;23;28m;[0m[38;2;84;84;91mh[0m[38;2;178;179;194m&[0m[38;2;187;188;205m&[0m[38;2;187;187;204m&[0m[38;2;188;189;205m&[0m[38;2;190;191;208m&[0m[38;2;194;194;212m&[0m[38;2;181;182;198m&[0m[38;2;72;74;81m3[0m[38;2;27;28;35mi[0m[38;2;22;24;30mi[0m[38;2;13;15;19m:[0m[38;2;4;5;7m.[0m[38;2;0;0;2m.[0m[38;2;24;24;25m;[0m[38;2;85;86;89mh[0m[38;2;149;150;154m9[0m[38;2;99;101;105mH[0m[38;2;0;0;0m [0m[38;2;10;10;11m,[0m[38;2;158;159;165m9[0m[38;2;243;246;252m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;244m@[0m");
    $display("[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;254;254;254m,[0m[38;2;170;170;170mi[0m[38;2;52;52;52m;[0m[38;2;2;2;2m,[0m[38;2;0;0;0m.[0m[38;2;1;2;3m.[0m[38;2;11;12;15m:[0m[38;2;19;20;25m;[0m[38;2;24;25;31mi[0m[38;2;27;28;35mi[0m[38;2;28;30;35mi[0m[38;2;17;17;18m:[0m[38;2;80;89;105mh[0m[38;2;131;148;174m9[0m[38;2;129;145;171m9[0m[38;2;130;146;171m9[0m[38;2;130;146;171m9[0m[38;2;132;148;174m9[0m[38;2;114;128;151mS[0m[38;2;39;43;49ms[0m[38;2;80;86;106mh[0m[38;2;128;143;169m9[0m[38;2;120;134;159m#[0m[38;2;113;127;149mS[0m[38;2;104;116;138mG[0m[38;2;91;102;120mH[0m[38;2;75;84;98mh[0m[38;2;55;62;73m2[0m[38;2;36;41;48ms[0m[38;2;22;24;29mi[0m[38;2;14;15;18m:[0m[38;2;16;16;18m:[0m[38;2;28;28;30mi[0m[38;2;48;48;53mX[0m[38;2;65;65;71m5[0m[38;2;76;76;83m3[0m[38;2;83;83;91mh[0m[38;2;85;85;93mh[0m[38;2;84;84;92mh[0m[38;2;83;83;91mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;91mh[0m[38;2;83;83;91mh[0m[38;2;84;84;93mh[0m[38;2;85;85;93mh[0m[38;2;82;82;90mh[0m[38;2;71;72;79m5[0m[38;2;50;50;55mA[0m[38;2;19;19;20m;[0m[38;2;1;1;1m.[0m[38;2;0;0;0m [0m[38;2;0;0;0m [0m[38;2;0;0;0m [0m[38;2;6;5;6m.[0m[38;2;19;19;21m;[0m[38;2;24;25;27mi[0m[38;2;28;29;31mi[0m[38;2;10;10;11m,[0m[38;2;0;0;0m [0m[38;2;12;13;15m:[0m[38;2;30;32;40mr[0m[38;2;39;40;46ms[0m[38;2;120;121;131mS[0m[38;2;186;187;204m&[0m[38;2;177;178;194m&[0m[38;2;163;163;177mB[0m[38;2;135;135;146m#[0m[38;2;113;113;122mG[0m[38;2;86;86;93mh[0m[38;2;26;27;29mi[0m[38;2;4;4;5m.[0m[38;2;20;20;21m;[0m[38;2;47;47;49mX[0m[38;2;94;94;96mM[0m[38;2;155;157;161m9[0m[38;2;187;189;195m&[0m[38;2;130;131;136mS[0m[38;2;48;48;51mX[0m[38;2;36;36;39mr[0m[38;2;64;64;67m2[0m[38;2;4;4;4m.[0m[38;2;56;56;59mA[0m[38;2;201;203;208m@[0m[38;2;243;246;251m@[0m[38;2;237;240;245m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m");
    $display("[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;216;216;216m;[0m[38;2;90;90;90mi[0m[38;2;4;4;4m,[0m[38;2;1;2;3m,[0m[38;2;16;17;21m:[0m[38;2;25;27;33mi[0m[38;2;29;31;39mr[0m[38;2;31;33;41mr[0m[38;2;31;33;41mr[0m[38;2;31;33;41mr[0m[38;2;30;32;39mr[0m[38;2;13;13;15m:[0m[38;2;22;24;29mi[0m[38;2;112;126;149mS[0m[38;2;128;143;169m9[0m[38;2;125;140;166m#[0m[38;2;124;139;165m#[0m[38;2;124;140;166m#[0m[38;2;118;133;157m#[0m[38;2;39;43;51ms[0m[38;2;2;2;3m.[0m[38;2;89;99;119mH[0m[38;2;126;142;169m#[0m[38;2;124;139;165m#[0m[38;2;124;140;166m#[0m[38;2;125;141;167m#[0m[38;2;126;142;168m#[0m[38;2;127;143;169m9[0m[38;2;126;142;168m#[0m[38;2;123;140;165m#[0m[38;2;117;132;157m#[0m[38;2;106;119;142mS[0m[38;2;88;99;118mH[0m[38;2;57;65;77m2[0m[38;2;7;8;9m,[0m[38;2;5;5;5m.[0m[38;2;14;14;15m:[0m[38;2;23;22;24m;[0m[38;2;43;42;46ms[0m[38;2;64;64;70m2[0m[38;2;79;79;86m3[0m[38;2;84;84;93mh[0m[38;2;84;84;93mh[0m[38;2;83;83;91mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;83;83;91mh[0m[38;2;85;85;93mh[0m[38;2;83;84;91mh[0m[38;2;62;62;69m2[0m[38;2;23;24;29mi[0m[38;2;8;9;11m,[0m[38;2;3;4;4m.[0m[38;2;1;1;1m.[0m[38;2;0;0;0m [0m[38;2;2;2;3m.[0m[38;2;2;2;3m.[0m[38;2;2;2;2m.[0m[38;2;5;5;5m.[0m[38;2;9;10;11m,[0m[38;2;11;12;17m:[0m[38;2;11;12;16m:[0m[38;2;6;7;11m,[0m[38;2;21;21;24m;[0m[38;2;49;49;54mX[0m[38;2;40;40;43ms[0m[38;2;38;38;40ms[0m[38;2;15;15;16m:[0m[38;2;7;6;6m,[0m[38;2;83;83;85mh[0m[38;2;133;134;138m#[0m[38;2;173;175;180mB[0m[38;2;204;206;211m@[0m[38;2;220;222;228m@[0m[38;2;219;221;227m@[0m[38;2;187;188;193m&[0m[38;2;128;128;132mS[0m[38;2;120;121;124mG[0m[38;2;164;166;170mB[0m[38;2;216;219;225m@[0m[38;2;148;149;156m9[0m[38;2;4;4;4m.[0m[38;2;0;0;0m [0m[38;2;31;31;32mr[0m[38;2;135;136;141m#[0m[38;2;228;231;236m@[0m[38;2;240;243;248m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m");
    $display("[38;2;253;253;253m.[0m[38;2;174;174;174mi[0m[38;2;35;35;35m;[0m[38;2;0;0;0m.[0m[38;2;17;18;22m;[0m[38;2;29;31;39mr[0m[38;2;31;33;41mr[0m[38;2;31;33;41mr[0m[38;2;30;32;40mr[0m[38;2;30;32;40mr[0m[38;2;30;32;40mr[0m[38;2;31;33;41mr[0m[38;2;20;22;26m;[0m[38;2;0;0;0m [0m[38;2;48;54;64mA[0m[38;2;126;143;168m#[0m[38;2;133;148;173m9[0m[38;2;133;148;171m9[0m[38;2;140;153;175m9[0m[38;2;155;166;186mB[0m[38;2;114;121;136mS[0m[38;2;4;4;5m.[0m[38;2;43;45;49mX[0m[38;2;174;181;193m&[0m[38;2;192;199;211m@[0m[38;2;192;198;209m&[0m[38;2;192;199;211m@[0m[38;2;192;198;210m&[0m[38;2;190;197;209m&[0m[38;2;187;193;206m&[0m[38;2;173;182;197m&[0m[38;2;159;169;187mB[0m[38;2;146;158;179mB[0m[38;2;137;151;174m9[0m[38;2;135;151;176m9[0m[38;2;98;111;133mG[0m[38;2;9;9;10m,[0m[38;2;39;43;49ms[0m[38;2;91;103;122mH[0m[38;2;63;72;86m5[0m[38;2;32;36;43mr[0m[38;2;11;13;15m:[0m[38;2;13;13;14m:[0m[38;2;32;32;35mr[0m[38;2;56;56;62mA[0m[38;2;74;75;82m3[0m[38;2;84;84;92mh[0m[38;2;85;85;93mh[0m[38;2;84;84;92mh[0m[38;2;84;84;92mh[0m[38;2;83;83;91mh[0m[38;2;83;83;91mh[0m[38;2;83;82;91mh[0m[38;2;83;83;91mh[0m[38;2;84;84;92mh[0m[38;2;83;83;91mh[0m[38;2;75;76;82m3[0m[38;2;59;60;67m2[0m[38;2;41;42;49ms[0m[38;2;31;33;41mr[0m[38;2;31;33;41mr[0m[38;2;30;32;40mr[0m[38;2;24;26;33mi[0m[38;2;18;18;23m;[0m[38;2;30;33;42mr[0m[38;2;38;43;53mX[0m[38;2;38;42;51ms[0m[38;2;9;10;12m,[0m[38;2;4;4;4m.[0m[38;2;31;32;34mr[0m[38;2;70;70;73m5[0m[38;2;93;93;96mM[0m[38;2;116;117;120mG[0m[38;2;141;142;146m#[0m[38;2;163;164;170mB[0m[38;2;191;193;198m&[0m[38;2;218;220;225m@[0m[38;2;112;113;116mG[0m[38;2;8;8;9m,[0m[38;2;162;163;169mB[0m[38;2;248;251;255m@[0m[38;2;241;244;249m@[0m[38;2;229;231;237m@[0m[38;2;217;220;226m@[0m[38;2;213;215;221m@[0m[38;2;219;221;226m@[0m[38;2;233;237;242m@[0m[38;2;243;246;251m@[0m[38;2;243;246;251m@[0m[38;2;241;245;249m@[0m[38;2;111;111;114mG[0m[38;2;0;0;0m [0m[38;2;2;2;3m.[0m[38;2;12;12;14m:[0m[38;2;7;7;9m,[0m[38;2;74;74;77m3[0m[38;2;204;207;213m@[0m[38;2;241;244;249m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m");
    $display("[38;2;167;167;167ms[0m[38;2;19;19;19m;[0m[38;2;0;0;0m [0m[38;2;19;20;23m;[0m[38;2;31;33;41mr[0m[38;2;30;32;40mr[0m[38;2;30;32;40mr[0m[38;2;30;32;40mr[0m[38;2;30;32;40mr[0m[38;2;30;32;40mr[0m[38;2;29;31;38mr[0m[38;2;26;27;34mi[0m[38;2;7;8;9m,[0m[38;2;0;0;0m [0m[38;2;80;85;94mh[0m[38;2;144;150;163m9[0m[38;2;165;169;179mB[0m[38;2;209;213;220m@[0m[38;2;230;233;238m@[0m[38;2;236;238;243m@[0m[38;2;115;115;120mG[0m[38;2;0;0;0m [0m[38;2;107;108;112mH[0m[38;2;238;240;245m@[0m[38;2;240;242;247m@[0m[38;2;239;242;246m@[0m[38;2;239;242;246m@[0m[38;2;239;242;246m@[0m[38;2;239;242;246m@[0m[38;2;239;242;246m@[0m[38;2;239;241;245m@[0m[38;2;236;239;243m@[0m[38;2;231;234;239m@[0m[38;2;222;226;232m@[0m[38;2;218;222;231m@[0m[38;2;124;128;137mS[0m[38;2;1;1;1m.[0m[38;2;75;80;88m3[0m[38;2;167;178;196m&[0m[38;2;157;168;189mB[0m[38;2;144;157;178m9[0m[38;2;119;131;150mS[0m[38;2;82;90;105mM[0m[38;2;42;47;55mX[0m[38;2;16;17;21m:[0m[38;2;8;8;10m,[0m[38;2;21;21;24m;[0m[38;2;41;42;46ms[0m[38;2;58;59;64m2[0m[38;2;67;68;75m5[0m[38;2;74;74;81m3[0m[38;2;77;77;85m3[0m[38;2;80;80;88m3[0m[38;2;76;75;83m3[0m[38;2;62;63;70m2[0m[38;2;48;48;56mX[0m[38;2;35;36;43ms[0m[38;2;29;31;39mr[0m[38;2;30;32;40mr[0m[38;2;31;33;41mr[0m[38;2;28;30;38mr[0m[38;2;25;26;33mi[0m[38;2;34;35;41mr[0m[38;2;88;95;108mM[0m[38;2;150;160;180mB[0m[38;2;174;184;200m&[0m[38;2;194;201;213m@[0m[38;2;104;105;111mH[0m[38;2;0;0;0m [0m[38;2;58;59;62m2[0m[38;2;213;216;222m@[0m[38;2;196;197;203m&[0m[38;2;149;151;157m9[0m[38;2;138;139;143m#[0m[38;2;134;134;134m#[0m[38;2;129;128;129mS[0m[38;2;126;126;128mS[0m[38;2;67;68;70m5[0m[38;2;0;0;0m [0m[38;2;85;85;88mh[0m[38;2;231;234;239m@[0m[38;2;236;239;244m@[0m[38;2;236;239;244m@[0m[38;2;237;240;244m@[0m[38;2;237;240;245m@[0m[38;2;237;240;245m@[0m[38;2;236;239;244m@[0m[38;2;235;238;243m@[0m[38;2;239;242;247m@[0m[38;2;219;221;226m@[0m[38;2;58;58;61m2[0m[38;2;0;0;0m [0m[38;2;16;16;17m:[0m[38;2;15;17;19m:[0m[38;2;67;77;89m3[0m[38;2;17;19;23m;[0m[38;2;41;41;43ms[0m[38;2;189;191;196m&[0m[38;2;241;244;249m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m");
    $display("[38;2;96;96;96mX[0m[38;2;0;0;0m.[0m[38;2;16;17;21m;[0m[38;2;32;34;42mr[0m[38;2;31;33;41mr[0m[38;2;31;33;41mr[0m[38;2;30;32;41mr[0m[38;2;30;32;40mr[0m[38;2;30;32;40mr[0m[38;2;30;32;40mr[0m[38;2;19;20;23m;[0m[38;2;2;3;3m.[0m[38;2;3;3;5m.[0m[38;2;7;10;17m,[0m[38;2;16;19;27m;[0m[38;2;12;13;15m:[0m[38;2;13;12;13m:[0m[38;2;128;128;131mS[0m[38;2;238;241;246m@[0m[38;2;230;233;238m@[0m[38;2;72;73;76m5[0m[38;2;2;2;2m.[0m[38;2;153;155;159m9[0m[38;2;241;244;249m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;236;239;244m@[0m[38;2;237;240;244m@[0m[38;2;244;247;251m@[0m[38;2;137;137;140m#[0m[38;2;0;0;0m [0m[38;2;111;109;111mH[0m[38;2;238;240;244m@[0m[38;2;235;238;243m@[0m[38;2;231;234;240m@[0m[38;2;227;230;237m@[0m[38;2;223;227;235m@[0m[38;2;211;216;225m@[0m[38;2;192;195;204m&[0m[38;2;156;159;165m9[0m[38;2;103;103;107mH[0m[38;2;48;48;50mX[0m[38;2;14;14;15m:[0m[38;2;4;4;5m.[0m[38;2;8;8;11m,[0m[38;2;19;20;24m;[0m[38;2;29;30;36mr[0m[38;2;31;32;39mr[0m[38;2;28;30;38mr[0m[38;2;28;30;38mr[0m[38;2;28;30;38mr[0m[38;2;25;26;33mi[0m[38;2;17;19;24m;[0m[38;2;10;11;15m:[0m[38;2;21;21;24m;[0m[38;2;93;93;96mM[0m[38;2;188;190;195m&[0m[38;2;227;231;238m@[0m[38;2;235;238;243m@[0m[38;2;239;241;245m@[0m[38;2;243;246;251m@[0m[38;2;194;196;201m&[0m[38;2;26;27;28mi[0m[38;2;5;5;6m.[0m[38;2;151;153;158m9[0m[38;2;127;127;132mS[0m[38;2;0;0;0m [0m[38;2;0;0;2m.[0m[38;2;14;22;47mi[0m[38;2;17;27;59mr[0m[38;2;11;17;36m;[0m[38;2;0;0;0m [0m[38;2;0;0;0m [0m[38;2;38;38;41ms[0m[38;2;208;210;216m@[0m[38;2;241;244;249m@[0m[38;2;238;241;246m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;236;239;244m@[0m[38;2;239;241;247m@[0m[38;2;128;129;133mS[0m[38;2;5;5;6m.[0m[38;2;24;24;26mi[0m[38;2;14;15;16m:[0m[38;2;8;8;8m,[0m[38;2;86;95;110mM[0m[38;2;110;124;146mS[0m[38;2;32;36;44mr[0m[38;2;38;37;38ms[0m[38;2;193;195;199m&[0m[38;2;241;244;249m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m");
    $display("[38;2;186;186;186mr[0m[38;2;42;42;42mi[0m[38;2;0;0;0m,[0m[38;2;8;9;13m:[0m[38;2;17;19;25mi[0m[38;2;21;22;29mi[0m[38;2;22;24;31mi[0m[38;2;25;27;34mi[0m[38;2;29;30;38mr[0m[38;2;28;30;38mr[0m[38;2;19;21;25m;[0m[38;2;0;0;0m [0m[38;2;12;16;26m:[0m[38;2;47;71;141mh[0m[38;2;48;73;147mh[0m[38;2;12;16;29m;[0m[38;2;3;2;1m.[0m[38;2;155;156;161m9[0m[38;2;249;252;255m@[0m[38;2;223;225;229m@[0m[38;2;49;49;50mX[0m[38;2;12;12;15m:[0m[38;2;175;175;180mB[0m[38;2;239;242;247m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;241;244;249m@[0m[38;2;141;141;145m#[0m[38;2;0;0;0m [0m[38;2;101;101;105mH[0m[38;2;240;242;247m@[0m[38;2;238;241;246m@[0m[38;2;236;239;244m@[0m[38;2;237;239;244m@[0m[38;2;237;240;245m@[0m[38;2;238;241;246m@[0m[38;2;240;243;248m@[0m[38;2;242;245;250m@[0m[38;2;242;245;250m@[0m[38;2;232;235;240m@[0m[38;2;204;206;211m@[0m[38;2;154;155;159m9[0m[38;2;99;100;103mM[0m[38;2;54;54;56mA[0m[38;2;25;25;27mi[0m[38;2;13;13;15m:[0m[38;2;7;8;9m,[0m[38;2;6;7;8m,[0m[38;2;6;7;8m,[0m[38;2;17;17;19m:[0m[38;2;44;45;46mX[0m[38;2;107;108;110mH[0m[38;2;188;190;194m&[0m[38;2;235;239;244m@[0m[38;2;241;244;249m@[0m[38;2;237;240;244m@[0m[38;2;236;238;243m@[0m[38;2;235;238;243m@[0m[38;2;237;240;244m@[0m[38;2;230;232;237m@[0m[38;2;78;79;82m3[0m[38;2;0;0;0m [0m[38;2;87;87;89mh[0m[38;2;145;146;152m9[0m[38;2;7;7;6m,[0m[38;2;8;11;16m,[0m[38;2;49;74;147mh[0m[38;2;57;89;183mH[0m[38;2;37;56;106m2[0m[38;2;0;0;0m [0m[38;2;0;0;0m [0m[38;2;13;12;12m:[0m[38;2;169;170;176mB[0m[38;2;224;226;232m@[0m[38;2;214;217;222m@[0m[38;2;233;236;241m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;237;240;245m@[0m[38;2;241;244;249m@[0m[38;2;156;157;161m9[0m[38;2;12;11;12m,[0m[38;2;50;51;54mA[0m[38;2;106;106;110mH[0m[38;2;6;6;6m,[0m[38;2;5;5;5m.[0m[38;2;73;81;95m3[0m[38;2;133;149;176m9[0m[38;2;123;138;163m#[0m[38;2;59;68;80m5[0m[38;2;57;58;61mA[0m[38;2;202;203;207m@[0m[38;2;240;243;248m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m");
    $display("[38;2;255;255;255m.[0m[38;2;224;224;224m:[0m[38;2;140;140;140mi[0m[38;2;80;79;79m;[0m[38;2;50;50;50m:[0m[38;2;38;38;38m:[0m[38;2;42;42;43m;[0m[38;2;34;34;35m;[0m[38;2;17;17;18m:[0m[38;2;55;55;56mr[0m[38;2;42;42;42mi[0m[38;2;0;0;0m [0m[38;2;22;31;56mr[0m[38;2;54;83;168mH[0m[38;2;54;83;170mH[0m[38;2;24;34;66ms[0m[38;2;4;4;4m.[0m[38;2;63;62;61m2[0m[38;2;111;111;111mH[0m[38;2;82;82;85m3[0m[38;2;10;10;10m,[0m[38;2;9;9;11m,[0m[38;2;160;162;166mB[0m[38;2;241;244;249m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;236;239;244m@[0m[38;2;237;240;245m@[0m[38;2;245;249;254m@[0m[38;2;138;139;142m#[0m[38;2;0;0;0m [0m[38;2;73;73;75m5[0m[38;2;189;190;196m&[0m[38;2;217;219;225m@[0m[38;2;236;239;244m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;238;241;246m@[0m[38;2;190;191;196m&[0m[38;2;141;142;147m#[0m[38;2;188;189;194m&[0m[38;2;223;226;232m@[0m[38;2;232;235;240m@[0m[38;2;222;225;230m@[0m[38;2;166;167;172mB[0m[38;2;23;22;23m;[0m[38;2;0;0;0m [0m[38;2;8;9;10m,[0m[38;2;146;148;153m9[0m[38;2;230;233;238m@[0m[38;2;241;244;249m@[0m[38;2;241;244;249m@[0m[38;2;236;239;244m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;237;240;245m@[0m[38;2;219;222;227m@[0m[38;2;68;69;72m5[0m[38;2;0;0;0m [0m[38;2;21;21;21m;[0m[38;2;39;39;39ms[0m[38;2;1;0;0m.[0m[38;2;30;42;79mX[0m[38;2;54;82;168mH[0m[38;2;55;86;175mH[0m[38;2;48;73;148mh[0m[38;2;21;31;59mr[0m[38;2;7;10;17m,[0m[38;2;3;3;4m.[0m[38;2;33;33;34mr[0m[38;2;36;36;38mr[0m[38;2;48;49;52mX[0m[38;2;200;203;208m@[0m[38;2;238;241;246m@[0m[38;2;239;242;247m@[0m[38;2;237;239;245m@[0m[38;2;144;145;150m9[0m[38;2;13;13;14m:[0m[38;2;38;38;40ms[0m[38;2;191;193;198m&[0m[38;2;139;140;144m#[0m[38;2;3;3;3m.[0m[38;2;9;9;9m,[0m[38;2;72;80;94m3[0m[38;2;130;146;172m9[0m[38;2;129;145;170m9[0m[38;2;129;145;171m9[0m[38;2;88;98;117mM[0m[38;2;91;93;101mM[0m[38;2;213;215;219m@[0m[38;2;239;242;247m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m");
    $display("[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m.[0m[38;2;248;248;248m,[0m[38;2;239;239;239m,[0m[38;2;239;239;239m:[0m[38;2;104;104;104ms[0m[38;2;2;2;2m.[0m[38;2;15;15;17m,[0m[38;2;14;16;23m:[0m[38;2;20;28;50mr[0m[38;2;48;71;142mh[0m[38;2;55;85;175mH[0m[38;2;54;84;173mH[0m[38;2;53;82;167mM[0m[38;2;44;67;134m3[0m[38;2;31;48;100m2[0m[38;2;22;35;75ms[0m[38;2;2;4;10m.[0m[38;2;0;0;0m [0m[38;2;0;0;0m [0m[38;2;85;86;89mh[0m[38;2;229;232;237m@[0m[38;2;237;240;245m@[0m[38;2;238;241;246m@[0m[38;2;239;242;247m@[0m[38;2;239;242;247m@[0m[38;2;241;245;250m@[0m[38;2;243;246;252m@[0m[38;2;243;246;251m@[0m[38;2;241;244;249m@[0m[38;2;235;238;243m@[0m[38;2;225;227;233m@[0m[38;2;199;201;206m@[0m[38;2;72;72;75m5[0m[38;2;0;0;0m [0m[38;2;6;6;6m,[0m[38;2;62;62;66m2[0m[38;2;203;206;212m@[0m[38;2;239;242;247m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;238;241;246m@[0m[38;2;197;199;205m&[0m[38;2;83;83;86mh[0m[38;2;38;38;39ms[0m[38;2;39;40;42ms[0m[38;2;67;68;71m5[0m[38;2;109;110;112mH[0m[38;2;115;116;121mG[0m[38;2;19;19;20m;[0m[38;2;2;3;3m.[0m[38;2;0;0;0m [0m[38;2;107;107;112mH[0m[38;2;237;240;246m@[0m[38;2;242;245;250m@[0m[38;2;243;246;251m@[0m[38;2;243;246;251m@[0m[38;2;242;245;250m@[0m[38;2;242;245;250m@[0m[38;2;240;243;248m@[0m[38;2;236;239;244m@[0m[38;2;240;243;248m@[0m[38;2;189;191;197m&[0m[38;2;18;18;20m;[0m[38;2;0;0;0m [0m[38;2;13;18;33m;[0m[38;2;20;29;58mr[0m[38;2;36;52;102m2[0m[38;2;54;83;170mH[0m[38;2;54;85;174mH[0m[38;2;54;84;172mH[0m[38;2;55;85;174mH[0m[38;2;55;86;176mH[0m[38;2;52;80;161mM[0m[38;2;47;72;145mh[0m[38;2;36;55;109m2[0m[38;2;2;5;11m,[0m[38;2;25;25;27mi[0m[38;2;190;192;196m&[0m[38;2;245;248;253m@[0m[38;2;222;225;231m@[0m[38;2;102;102;105mH[0m[38;2;4;4;5m.[0m[38;2;66;66;69m5[0m[38;2;200;202;208m@[0m[38;2;241;244;250m@[0m[38;2;99;100;106mH[0m[38;2;1;1;1m [0m[38;2;26;26;26m;[0m[38;2;80;89;103mh[0m[38;2;129;146;171m9[0m[38;2;127;143;168m#[0m[38;2;127;143;168m#[0m[38;2;130;147;173m9[0m[38;2;111;124;147mS[0m[38;2;125;130;141mS[0m[38;2;221;223;228m@[0m[38;2;238;241;245m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m");
    $display("[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m.[0m[38;2;111;111;111ms[0m[38;2;0;0;0m.[0m[38;2;14;20;39mi[0m[38;2;32;49;99m2[0m[38;2;42;63;124m3[0m[38;2;53;82;166mM[0m[38;2;54;85;174mH[0m[38;2;54;84;172mH[0m[38;2;55;85;174mH[0m[38;2;53;81;165mM[0m[38;2;47;72;147mh[0m[38;2;39;59;118m5[0m[38;2;12;16;28m;[0m[38;2;0;0;0m [0m[38;2;0;0;1m.[0m[38;2;8;8;10m,[0m[38;2;160;162;167mB[0m[38;2;243;245;251m@[0m[38;2;213;215;220m@[0m[38;2;207;210;214m@[0m[38;2;204;206;211m@[0m[38;2;170;172;176mB[0m[38;2;132;134;139m#[0m[38;2;106;108;111mH[0m[38;2;85;86;89mh[0m[38;2;63;64;66m2[0m[38;2;44;44;47mX[0m[38;2;29;30;31mi[0m[38;2;3;3;4m.[0m[38;2;0;0;0m [0m[38;2;0;1;2m.[0m[38;2;138;139;144m#[0m[38;2;241;244;249m@[0m[38;2;233;236;241m@[0m[38;2;237;240;245m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;238;242;247m@[0m[38;2;238;241;246m@[0m[38;2;217;220;224m@[0m[38;2;182;184;189m&[0m[38;2;140;141;146m#[0m[38;2;100;101;104mH[0m[38;2;57;58;60mA[0m[38;2;6;7;7m,[0m[38;2;10;8;8m,[0m[38;2;5;4;4m.[0m[38;2;14;14;15m:[0m[38;2;70;70;74m5[0m[38;2;98;98;102mM[0m[38;2;119;121;125mG[0m[38;2;140;142;146m#[0m[38;2;158;160;165mB[0m[38;2;171;173;178mB[0m[38;2;189;191;195m&[0m[38;2;226;228;233m@[0m[38;2;243;246;252m@[0m[38;2;218;220;226m@[0m[38;2;60;60;61m2[0m[38;2;0;0;0m [0m[38;2;16;23;40mi[0m[38;2;18;29;60mr[0m[38;2;26;38;74mX[0m[38;2;43;64;128m3[0m[38;2;54;84;172mH[0m[38;2;54;85;174mH[0m[38;2;54;84;173mH[0m[38;2;48;73;146mh[0m[38;2;38;57;112m5[0m[38;2;31;45;87mA[0m[38;2;26;37;70ms[0m[38;2;2;4;10m.[0m[38;2;9;9;9m,[0m[38;2;180;182;187m&[0m[38;2;205;207;213m@[0m[38;2;62;62;66m2[0m[38;2;15;15;16m:[0m[38;2;122;123;127mS[0m[38;2;224;227;232m@[0m[38;2;241;244;249m@[0m[38;2;234;237;243m@[0m[38;2;83;84;87mh[0m[38;2;0;0;0m [0m[38;2;30;32;36mr[0m[38;2;101;113;134mG[0m[38;2;129;145;171m9[0m[38;2;127;143;168m#[0m[38;2;127;143;168m#[0m[38;2;127;143;168m#[0m[38;2;129;145;170m9[0m[38;2;117;132;156m#[0m[38;2;141;146;159m9[0m[38;2;225;228;233m@[0m[38;2;237;240;245m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m");
    $display("[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;209;209;209m;[0m[38;2;77;77;77mi[0m[38;2;34;34;35m;[0m[38;2;40;40;41m;[0m[38;2;6;6;6m.[0m[38;2;19;26;49mr[0m[38;2;52;79;160mM[0m[38;2;57;89;183mH[0m[38;2;42;61;121m5[0m[38;2;10;13;24m:[0m[38;2;9;9;12m,[0m[38;2;29;30;31mi[0m[38;2;24;25;27mi[0m[38;2;9;9;10m,[0m[38;2;3;3;4m.[0m[38;2;19;16;16m:[0m[38;2;53;54;56mA[0m[38;2;172;173;178mB[0m[38;2;55;55;57mA[0m[38;2;49;50;53mX[0m[38;2;105;105;109mH[0m[38;2;97;97;100mM[0m[38;2;96;98;102mM[0m[38;2;109;110;113mH[0m[38;2;131;133;137m#[0m[38;2;155;157;161m9[0m[38;2;184;186;191m&[0m[38;2;195;197;202m&[0m[38;2;57;57;60mA[0m[38;2;23;22;24m;[0m[38;2;12;11;12m,[0m[38;2;62;63;66m2[0m[38;2;191;192;198m&[0m[38;2;85;86;90mh[0m[38;2;181;185;190m&[0m[38;2;246;249;255m@[0m[38;2;243;246;251m@[0m[38;2;243;246;251m@[0m[38;2;242;245;251m@[0m[38;2;242;245;250m@[0m[38;2;241;244;250m@[0m[38;2;241;244;249m@[0m[38;2;242;245;250m@[0m[38;2;244;246;252m@[0m[38;2;245;248;254m@[0m[38;2;251;255;255m@[0m[38;2;178;181;187m&[0m[38;2;17;20;23m;[0m[38;2;131;94;91mH[0m[38;2;148;106;98mG[0m[38;2;65;64;68m2[0m[38;2;163;165;171mB[0m[38;2;151;151;155m9[0m[38;2;132;133;138m#[0m[38;2;124;125;130mS[0m[38;2;121;122;127mS[0m[38;2;127;128;133mS[0m[38;2;154;154;160m9[0m[38;2;190;192;196m&[0m[38;2;201;203;207m@[0m[38;2;201;203;207m@[0m[38;2;153;156;160m9[0m[38;2;16;16;16m:[0m[38;2;6;6;5m.[0m[38;2;76;75;74m3[0m[38;2;21;19;17m;[0m[38;2;4;5;7m.[0m[38;2;41;60;116m5[0m[38;2;54;84;172mH[0m[38;2;51;77;155mM[0m[38;2;18;23;40mi[0m[38;2;0;0;0m [0m[38;2;0;0;0m [0m[38;2;6;5;3m.[0m[38;2;65;65;67m2[0m[38;2;99;99;103mM[0m[38;2;112;113;119mG[0m[38;2;45;46;49mX[0m[38;2;77;78;82m3[0m[38;2;191;193;198m&[0m[38;2;240;243;248m@[0m[38;2;238;241;246m@[0m[38;2;238;241;246m@[0m[38;2;215;217;223m@[0m[38;2;49;49;52mX[0m[38;2;0;0;0m [0m[38;2;17;18;21m;[0m[38;2;109;123;145mS[0m[38;2;129;145;171m9[0m[38;2;127;143;168m#[0m[38;2;127;143;168m#[0m[38;2;127;143;168m#[0m[38;2;127;143;168m#[0m[38;2;128;144;169m9[0m[38;2;117;132;157m#[0m[38;2;158;166;182mB[0m[38;2;233;236;241m@[0m[38;2;236;239;244m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m");
    $display("[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;251;251;250m,[0m[38;2;234;234;234m:[0m[38;2;212;212;212mi[0m[38;2;32;31;31m;[0m[38;2;0;0;0m [0m[38;2;19;29;58mr[0m[38;2;22;37;78mX[0m[38;2;9;14;32m;[0m[38;2;0;0;0m [0m[38;2;12;12;12m:[0m[38;2;155;156;162m9[0m[38;2;214;217;223m@[0m[38;2;84;84;89mh[0m[38;2;0;0;0m [0m[38;2;72;57;56m2[0m[38;2;124;96;92mH[0m[38;2;51;49;52mX[0m[38;2;15;13;15m:[0m[38;2;27;28;31mi[0m[38;2;153;155;159m9[0m[38;2;178;180;184m&[0m[38;2;172;174;179mB[0m[38;2;170;172;177mB[0m[38;2;168;170;175mB[0m[38;2;163;165;170mB[0m[38;2;161;163;169mB[0m[38;2;172;174;179mB[0m[38;2;96;98;103mM[0m[38;2;123;114;112mG[0m[38;2;170;157;151m9[0m[38;2;46;44;45mX[0m[38;2;64;65;69m2[0m[38;2;52;40;40ms[0m[38;2;127;114;115mG[0m[38;2;122;123;128mS[0m[38;2;103;106;110mH[0m[38;2;99;101;105mH[0m[38;2;94;96;100mM[0m[38;2;88;90;95mh[0m[38;2;84;85;89mh[0m[38;2;84;85;88mh[0m[38;2;81;81;84m3[0m[38;2;81;80;83m3[0m[38;2;91;89;90mh[0m[38;2;119;115;117mG[0m[38;2;95;89;92mM[0m[38;2;102;77;73mh[0m[38;2;241;188;175m@[0m[38;2;255;209;194m@[0m[38;2;152;129;126m#[0m[38;2;71;71;73m5[0m[38;2;51;51;52mX[0m[38;2;52;50;51mX[0m[38;2;54;52;54mA[0m[38;2;49;48;50mX[0m[38;2;44;45;47mX[0m[38;2;37;37;39ms[0m[38;2;18;18;18m:[0m[38;2;11;11;11m,[0m[38;2;22;21;22m;[0m[38;2;60;52;52mA[0m[38;2;13;10;11m,[0m[38;2;20;20;21m;[0m[38;2;163;163;169mB[0m[38;2;53;53;57mA[0m[38;2;0;0;0m [0m[38;2;5;7;14m,[0m[38;2;10;15;31m;[0m[38;2;7;11;24m:[0m[38;2;4;4;6m.[0m[38;2;20;21;22m;[0m[38;2;8;9;9m,[0m[38;2;25;25;27mi[0m[38;2;166;167;173mB[0m[38;2;129;130;135mS[0m[38;2;101;102;106mH[0m[38;2;180;182;187m&[0m[38;2;237;239;245m@[0m[38;2;240;243;248m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;241;244;249m@[0m[38;2;146;147;151m9[0m[38;2;5;5;5m,[0m[38;2;6;6;6m,[0m[38;2;3;3;3m.[0m[38;2;72;82;96mh[0m[38;2;128;145;170m9[0m[38;2;127;143;168m#[0m[38;2;127;143;168m#[0m[38;2;127;143;168m#[0m[38;2;127;143;168m#[0m[38;2;127;143;168m#[0m[38;2;127;143;168m#[0m[38;2;125;140;164m#[0m[38;2;186;192;204m&[0m[38;2;237;240;244m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m");
    $display("[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;236;236;236m:[0m[38;2;57;57;57mr[0m[38;2;0;0;0m [0m[38;2;44;43;44ms[0m[38;2;75;75;75m3[0m[38;2;83;83;85mh[0m[38;2;130;131;135mS[0m[38;2;183;185;190m&[0m[38;2;227;230;235m@[0m[38;2;244;247;252m@[0m[38;2;129;129;132mS[0m[38;2;0;0;0m [0m[38;2;37;28;28mr[0m[38;2;206;151;142mB[0m[38;2;147;116;110mS[0m[38;2;159;126;120m#[0m[38;2;139;112;107mG[0m[38;2;89;79;77m3[0m[38;2;73;69;67m5[0m[38;2;70;65;64m2[0m[38;2;69;65;63m2[0m[38;2;69;64;63m2[0m[38;2;69;65;63m2[0m[38;2;70;65;63m2[0m[38;2;82;77;75m3[0m[38;2;120;113;110mG[0m[38;2;165;154;149m9[0m[38;2;173;162;156mB[0m[38;2;94;88;87mh[0m[38;2;13;14;17m:[0m[38;2;144;111;105mG[0m[38;2;220;175;164m&[0m[38;2;109;93;89mM[0m[38;2;113;91;88mM[0m[38;2;120;100;96mH[0m[38;2;122;103;98mH[0m[38;2;133;110;104mG[0m[38;2;126;102;97mH[0m[38;2;24;20;20m;[0m[38;2;0;0;0m [0m[38;2;13;9;10m,[0m[38;2;59;44;43mX[0m[38;2;95;68;64m3[0m[38;2;113;92;88mM[0m[38;2;146;125;121mS[0m[38;2;149;138;133m#[0m[38;2;147;138;133m#[0m[38;2;130;119;114mG[0m[38;2;73;68;67m5[0m[38;2;33;32;35mr[0m[38;2;30;24;27mi[0m[38;2;29;23;24mi[0m[38;2;11;9;12m,[0m[38;2;0;0;1m.[0m[38;2;0;0;0m [0m[38;2;0;0;0m [0m[38;2;0;0;0m [0m[38;2;62;52;53mA[0m[38;2;188;138;129m9[0m[38;2;37;26;23mi[0m[38;2;16;17;19m:[0m[38;2;170;171;176mB[0m[38;2;176;177;182m&[0m[38;2;157;158;164m9[0m[38;2;153;155;159m9[0m[38;2;150;151;152m9[0m[38;2;150;151;154m9[0m[38;2;172;173;178mB[0m[38;2;196;198;203m&[0m[38;2;56;56;59mA[0m[38;2;5;5;5m.[0m[38;2;105;105;109mH[0m[38;2;205;207;212m@[0m[38;2;239;242;247m@[0m[38;2;241;244;249m@[0m[38;2;236;239;244m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;241;244;249m@[0m[38;2;203;206;211m@[0m[38;2;40;40;43ms[0m[38;2;25;25;25m:[0m[38;2;119;119;119mX[0m[38;2;15;15;15m,[0m[38;2;26;29;35mr[0m[38;2;116;130;154mS[0m[38;2;128;145;170m9[0m[38;2;127;143;168m#[0m[38;2;127;143;168m#[0m[38;2;127;143;168m#[0m[38;2;127;143;168m#[0m[38;2;127;143;168m#[0m[38;2;126;142;168m#[0m[38;2;135;148;170m9[0m[38;2;206;209;218m@[0m[38;2;238;240;245m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m");
    $display("[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;248;248;248m:[0m[38;2;87;87;87ms[0m[38;2;0;0;0m.[0m[38;2;143;144;151m#[0m[38;2;242;245;251m@[0m[38;2;240;243;248m@[0m[38;2;242;246;251m@[0m[38;2;241;244;249m@[0m[38;2;236;239;244m@[0m[38;2;240;243;248m@[0m[38;2;183;185;190m&[0m[38;2;18;18;19m;[0m[38;2;2;1;1m.[0m[38;2;32;28;28mi[0m[38;2;27;24;24mi[0m[38;2;35;33;32mr[0m[38;2;55;50;49mX[0m[38;2;60;55;53mA[0m[38;2;61;58;56mA[0m[38;2;67;64;63m2[0m[38;2;72;69;68m5[0m[38;2;67;64;63m2[0m[38;2;58;54;55mA[0m[38;2;50;46;47mX[0m[38;2;38;35;36mr[0m[38;2;26;23;25mi[0m[38;2;7;6;9m,[0m[38;2;0;0;0m [0m[38;2;0;0;0m [0m[38;2;2;3;4m.[0m[38;2;156;146;141m9[0m[38;2;255;241;229m@[0m[38;2;255;240;229m@[0m[38;2;255;241;230m@[0m[38;2;255;242;230m@[0m[38;2;255;242;230m@[0m[38;2;255;242;231m@[0m[38;2;255;238;227m@[0m[38;2;199;185;176m&[0m[38;2;141;131;127mS[0m[38;2;107;100;96mM[0m[38;2;82;78;76m3[0m[38;2;69;65;64m2[0m[38;2;54;52;50mA[0m[38;2;43;43;44ms[0m[38;2;40;40;40ms[0m[38;2;17;18;19m:[0m[38;2;0;0;0m [0m[38;2;15;15;15m:[0m[38;2;48;50;37ms[0m[38;2;51;52;40mX[0m[38;2;62;65;48mA[0m[38;2;77;80;53m5[0m[38;2;98;101;69mh[0m[38;2;116;120;83mH[0m[38;2;36;36;31mr[0m[38;2;1;2;4m.[0m[38;2;164;151;147m9[0m[38;2;224;190;179m&[0m[38;2;30;22;21m;[0m[38;2;21;22;24m;[0m[38;2;192;194;198m&[0m[38;2;246;249;254m@[0m[38;2;242;246;251m@[0m[38;2;243;246;251m@[0m[38;2;243;246;251m@[0m[38;2;243;246;251m@[0m[38;2;243;247;251m@[0m[38;2;229;232;237m@[0m[38;2;70;70;72m5[0m[38;2;0;0;0m [0m[38;2;42;42;44ms[0m[38;2;178;181;186m&[0m[38;2;240;243;248m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;240;244;249m@[0m[38;2;217;218;223m@[0m[38;2;73;73;75m5[0m[38;2;3;3;3m,[0m[38;2;147;147;147mr[0m[38;2;242;242;242m;[0m[38;2;72;71;72mr[0m[38;2;0;0;0m.[0m[38;2;81;91;108mM[0m[38;2;130;146;171m9[0m[38;2;127;143;168m#[0m[38;2;127;143;168m#[0m[38;2;127;143;168m#[0m[38;2;127;143;168m#[0m[38;2;127;143;168m#[0m[38;2;127;143;168m#[0m[38;2;125;141;166m#[0m[38;2;144;156;176m9[0m[38;2;217;221;227m@[0m[38;2;237;240;245m@[0m[38;2;235;238;243m@[0m");
    $display("[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;246;246;246m:[0m[38;2;85;85;86ms[0m[38;2;0;0;0m.[0m[38;2;141;143;149m#[0m[38;2;240;243;248m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;236;239;244m@[0m[38;2;231;234;239m@[0m[38;2;95;95;99mM[0m[38;2;0;0;0m [0m[38;2;69;66;65m2[0m[38;2;158;147;142m9[0m[38;2;116;109;106mH[0m[38;2;85;80;78m3[0m[38;2;67;64;63m2[0m[38;2;62;59;58m2[0m[38;2;32;31;31mr[0m[38;2;0;0;0m [0m[38;2;13;14;12m,[0m[38;2;60;62;42mA[0m[38;2;69;72;48m2[0m[38;2;83;86;60m3[0m[38;2;100;104;71mh[0m[38;2;126;130;91mG[0m[38;2;129;135;94mG[0m[38;2;25;26;25mi[0m[38;2;11;12;13m:[0m[38;2;190;178;172m&[0m[38;2;255;240;228m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;254;236;225m@[0m[38;2;255;240;229m@[0m[38;2;255;243;232m@[0m[38;2;255;242;231m@[0m[38;2;255;240;229m@[0m[38;2;255;237;226m@[0m[38;2;249;231;220m@[0m[38;2;245;228;219m@[0m[38;2;247;232;221m@[0m[38;2;193;181;175m&[0m[38;2;25;25;27mi[0m[38;2;22;23;21m;[0m[38;2;157;162;113m#[0m[38;2;211;220;143m&[0m[38;2;212;221;143m&[0m[38;2;212;222;142m&[0m[38;2;220;229;147m&[0m[38;2;150;156;107m#[0m[38;2;10;10;9m,[0m[38;2;39;38;40ms[0m[38;2;222;206;197m@[0m[38;2;205;186;177m&[0m[38;2;19;14;13m:[0m[38;2;32;33;35mr[0m[38;2;200;202;207m@[0m[38;2;239;242;247m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;236;239;244m@[0m[38;2;231;234;239m@[0m[38;2;81;81;84m3[0m[38;2;0;0;1m.[0m[38;2;0;0;0m [0m[38;2;31;31;33mr[0m[38;2;186;188;193m&[0m[38;2;239;242;247m@[0m[38;2;235;238;243m@[0m[38;2;242;245;250m@[0m[38;2;208;210;215m@[0m[38;2;67;67;71m5[0m[38;2;2;2;1m,[0m[38;2;128;128;128mr[0m[38;2;251;251;251m,[0m[38;2;255;255;255m [0m[38;2;158;158;158ms[0m[38;2;5;5;4m,[0m[38;2;38;43;51ms[0m[38;2;122;138;162m#[0m[38;2;128;144;169m9[0m[38;2;127;143;168m#[0m[38;2;127;143;168m#[0m[38;2;127;143;168m#[0m[38;2;127;143;168m#[0m[38;2;127;143;168m#[0m[38;2;127;143;168m#[0m[38;2;124;140;166m#[0m[38;2;158;168;186mB[0m[38;2;230;232;237m@[0m[38;2;236;239;244m@[0m");
    $display("[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;250;250;250m,[0m[38;2;97;97;97ms[0m[38;2;0;0;0m.[0m[38;2;133;135;141m#[0m[38;2;239;241;247m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;240;243;248m@[0m[38;2;194;196;201m&[0m[38;2;31;31;33mr[0m[38;2;21;20;20m;[0m[38;2;205;190;183m&[0m[38;2;255;248;237m@[0m[38;2;255;240;229m@[0m[38;2;255;237;226m@[0m[38;2;255;239;228m@[0m[38;2;216;202;194m@[0m[38;2;52;49;50mX[0m[38;2;10;10;10m,[0m[38;2;126;131;92mG[0m[38;2;209;218;142m&[0m[38;2;218;227;146m&[0m[38;2;217;227;145m&[0m[38;2;216;225;145m&[0m[38;2;112;117;81mH[0m[38;2;0;0;0m [0m[38;2;78;74;73m3[0m[38;2;240;223;212m@[0m[38;2;254;237;226m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;254;236;225m@[0m[38;2;254;236;225m@[0m[38;2;255;237;225m@[0m[38;2;255;237;226m@[0m[38;2;255;239;227m@[0m[38;2;174;164;159mB[0m[38;2;32;30;31mr[0m[38;2;20;21;17m;[0m[38;2;106;111;78mM[0m[38;2;166;173;115m9[0m[38;2;181;189;123mB[0m[38;2;128;134;89mG[0m[38;2;20;22;17m;[0m[38;2;25;24;26mi[0m[38;2;172;162;158mB[0m[38;2;255;243;231m@[0m[38;2;169;158;152m9[0m[38;2;5;4;5m.[0m[38;2;52;52;56mA[0m[38;2;215;218;224m@[0m[38;2;238;241;246m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;236;239;244m@[0m[38;2;231;234;239m@[0m[38;2;79;78;81m3[0m[38;2;7;6;8m,[0m[38;2;54;54;58mA[0m[38;2;0;1;1m.[0m[38;2;82;83;86mh[0m[38;2;228;231;236m@[0m[38;2;244;247;253m@[0m[38;2;183;184;189m&[0m[38;2;42;42;45mX[0m[38;2;13;12;12m,[0m[38;2;140;140;140mr[0m[38;2;250;250;250m,[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;223;223;223mi[0m[38;2;46;45;45mi[0m[38;2;7;8;11m,[0m[38;2;99;112;132mG[0m[38;2;130;146;172m9[0m[38;2;127;143;168m#[0m[38;2;127;143;168m#[0m[38;2;127;143;168m#[0m[38;2;127;143;168m#[0m[38;2;127;143;168m#[0m[38;2;127;143;168m#[0m[38;2;127;143;168m#[0m[38;2;126;142;167m#[0m[38;2;187;193;205m&[0m[38;2;237;239;244m@[0m");
    $display("[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;254;254;254m.[0m[38;2;113;113;113ms[0m[38;2;0;0;0m.[0m[38;2;124;125;131mS[0m[38;2;245;248;254m@[0m[38;2;244;247;252m@[0m[38;2;243;246;251m@[0m[38;2;242;245;250m@[0m[38;2;240;243;248m@[0m[38;2;238;241;246m@[0m[38;2;237;240;245m@[0m[38;2;239;242;247m@[0m[38;2;134;135;139m#[0m[38;2;0;1;1m.[0m[38;2;83;78;76m3[0m[38;2;244;227;217m@[0m[38;2;255;237;226m@[0m[38;2;254;236;225m@[0m[38;2;254;236;225m@[0m[38;2;255;240;228m@[0m[38;2;217;202;194m@[0m[38;2;78;73;72m5[0m[38;2;8;8;10m,[0m[38;2;63;65;49mA[0m[38;2;140;145;99mS[0m[38;2;154;158;111m#[0m[38;2;84;88;61m3[0m[38;2;4;5;5m.[0m[38;2;64;61;61m2[0m[38;2;214;199;191m@[0m[38;2;255;239;228m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;254;236;225m@[0m[38;2;255;240;229m@[0m[38;2;222;206;197m@[0m[38;2;127;119;116mG[0m[38;2;56;53;55mA[0m[38;2;40;38;38mr[0m[38;2;41;41;38ms[0m[38;2;43;42;42ms[0m[38;2;102;96;94mM[0m[38;2;208;194;186m&[0m[38;2;255;239;228m@[0m[38;2;255;241;230m@[0m[38;2;155;143;139m#[0m[38;2;1;1;1m.[0m[38;2;81;81;84m3[0m[38;2;231;234;239m@[0m[38;2;236;239;244m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;236;240;245m@[0m[38;2;229;231;236m@[0m[38;2;70;70;72m5[0m[38;2;11;10;11m,[0m[38;2;137;129;127mS[0m[38;2;37;35;35mr[0m[38;2;21;21;22m;[0m[38;2;183;185;190m&[0m[38;2;140;142;146m9[0m[38;2;22;22;23mi[0m[38;2;69;69;69m;[0m[38;2;196;196;196mi[0m[38;2;255;255;255m.[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;254;254;254m.[0m[38;2;116;116;116ms[0m[38;2;0;0;0m.[0m[38;2;64;71;84m5[0m[38;2;128;144;170m9[0m[38;2;127;143;168m#[0m[38;2;127;143;168m#[0m[38;2;127;143;168m#[0m[38;2;127;143;168m#[0m[38;2;127;143;168m#[0m[38;2;127;143;168m#[0m[38;2;127;143;168m#[0m[38;2;125;142;167m#[0m[38;2;138;151;173m9[0m[38;2;211;214;222m@[0m");
    $display("[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m.[0m[38;2;135;135;134ms[0m[38;2;0;0;0m.[0m[38;2;89;90;95mh[0m[38;2;135;135;141m#[0m[38;2;107;108;112mH[0m[38;2;132;134;138m#[0m[38;2;167;169;174mB[0m[38;2;197;199;204m&[0m[38;2;218;221;226m@[0m[38;2;232;235;240m@[0m[38;2;242;245;251m@[0m[38;2;226;228;234m@[0m[38;2;65;66;69m2[0m[38;2;5;5;6m.[0m[38;2;170;159;154mB[0m[38;2;255;244;233m@[0m[38;2;255;237;226m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;255;240;228m@[0m[38;2;248;231;220m@[0m[38;2;173;162;157mB[0m[38;2;87;82;82mh[0m[38;2;49;46;48mX[0m[38;2;44;41;43ms[0m[38;2;66;61;62m2[0m[38;2;148;138;134m#[0m[38;2;238;221;211m@[0m[38;2;255;239;228m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;255;237;226m@[0m[38;2;255;241;229m@[0m[38;2;255;237;226m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;255;239;228m@[0m[38;2;255;242;231m@[0m[38;2;248;231;221m@[0m[38;2;230;214;205m@[0m[38;2;220;200;192m@[0m[38;2;237;214;205m@[0m[38;2;255;241;230m@[0m[38;2;255;240;228m@[0m[38;2;254;236;225m@[0m[38;2;254;237;226m@[0m[38;2;121;109;105mG[0m[38;2;0;0;0m [0m[38;2;114;115;120mG[0m[38;2;236;239;245m@[0m[38;2;236;239;244m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;237;240;245m@[0m[38;2;219;221;227m@[0m[38;2;54;54;57mA[0m[38;2;18;18;18m:[0m[38;2;164;152;146m9[0m[38;2;45;41;41ms[0m[38;2;1;2;3m,[0m[38;2;53;54;57m2[0m[38;2;59;59;59mi[0m[38;2;161;161;161m;[0m[38;2;248;248;248m,[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;184;184;184mr[0m[38;2;13;12;12m:[0m[38;2;30;33;39mr[0m[38;2;119;134;158m#[0m[38;2;128;144;170m9[0m[38;2;127;143;168m#[0m[38;2;127;143;168m#[0m[38;2;127;143;168m#[0m[38;2;127;143;168m#[0m[38;2;127;143;168m#[0m[38;2;127;143;168m#[0m[38;2;127;143;168m#[0m[38;2;125;141;167m#[0m[38;2;159;168;185mB[0m");
    $display("[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;164;164;164ms[0m[38;2;9;9;9m:[0m[38;2;25;25;27mi[0m[38;2;2;2;3m.[0m[38;2;25;24;25mi[0m[38;2;73;69;67m5[0m[38;2;53;50;50mX[0m[38;2;42;41;42ms[0m[38;2;44;44;46mX[0m[38;2;56;57;60mA[0m[38;2;76;77;81m3[0m[38;2;104;105;108mH[0m[38;2;72;73;77m5[0m[38;2;0;0;2m.[0m[38;2;51;48;49mX[0m[38;2;195;182;175m&[0m[38;2;250;232;222m@[0m[38;2;255;243;231m@[0m[38;2;255;238;227m@[0m[38;2;253;235;224m@[0m[38;2;255;236;225m@[0m[38;2;255;242;230m@[0m[38;2;255;239;228m@[0m[38;2;244;226;217m@[0m[38;2;238;222;212m@[0m[38;2;252;234;223m@[0m[38;2;255;242;231m@[0m[38;2;255;238;226m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;254;236;225m@[0m[38;2;233;217;207m@[0m[38;2;188;175;169mB[0m[38;2;232;215;205m@[0m[38;2;254;237;225m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;254;236;225m@[0m[38;2;255;239;228m@[0m[38;2;255;242;230m@[0m[38;2;255;240;229m@[0m[38;2;254;236;225m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;255;237;226m@[0m[38;2;255;237;226m@[0m[38;2;228;149;150mB[0m[38;2;220;126;130m9[0m[38;2;251;223;214m@[0m[38;2;253;237;225m@[0m[38;2;255;237;226m@[0m[38;2;243;225;215m@[0m[38;2;70;65;65m2[0m[38;2;3;4;4m.[0m[38;2;160;160;165mB[0m[38;2;241;243;249m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;239;242;247m@[0m[38;2;201;203;209m@[0m[38;2;35;35;37mr[0m[38;2;12;12;12m,[0m[38;2;44;43;44ms[0m[38;2;8;8;8m:[0m[38;2;71;71;72m;[0m[38;2;173;173;173m;[0m[38;2;243;243;243m,[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;231;231;231m;[0m[38;2;50;50;50mr[0m[38;2;8;8;11m,[0m[38;2;100;113;133mG[0m[38;2;130;146;171m9[0m[38;2;127;143;168m#[0m[38;2;127;143;168m#[0m[38;2;127;143;168m#[0m[38;2;127;143;168m#[0m[38;2;127;143;168m#[0m[38;2;127;143;168m#[0m[38;2;127;143;168m#[0m[38;2;127;143;168m#[0m[38;2;130;144;169m9[0m");
    $display("[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;205;205;205mi[0m[38;2;27;27;27m;[0m[38;2;5;5;6m,[0m[38;2;0;0;0m [0m[38;2;82;80;82m3[0m[38;2;246;230;221m@[0m[38;2;248;230;220m@[0m[38;2;229;213;204m@[0m[38;2;205;191;182m&[0m[38;2;179;166;160mB[0m[38;2;149;138;133m#[0m[38;2;132;124;120mS[0m[38;2;133;124;119mS[0m[38;2;168;158;154m9[0m[38;2;115;109;106mH[0m[38;2;34;32;33mr[0m[38;2;67;64;62m2[0m[38;2;155;145;141m9[0m[38;2;235;218;209m@[0m[38;2;255;239;228m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;254;236;225m@[0m[38;2;255;237;226m@[0m[38;2;255;237;226m@[0m[38;2;254;236;225m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;254;237;226m@[0m[38;2;209;194;186m&[0m[38;2;142;132;129m#[0m[38;2;225;209;200m@[0m[38;2;254;237;226m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;254;236;225m@[0m[38;2;255;239;227m@[0m[38;2;255;243;231m@[0m[38;2;255;237;226m@[0m[38;2;217;203;194m@[0m[38;2;181;169;162mB[0m[38;2;204;189;181m&[0m[38;2;250;231;221m@[0m[38;2;253;236;225m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;253;236;225m@[0m[38;2;251;228;217m@[0m[38;2;219;133;133mB[0m[38;2;212;108;114m#[0m[38;2;246;208;200m@[0m[38;2;254;238;226m@[0m[38;2;255;239;228m@[0m[38;2;212;195;186m&[0m[38;2;28;24;24mi[0m[38;2;30;30;31mi[0m[38;2;199;201;207m@[0m[38;2;239;242;247m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;240;244;249m@[0m[38;2;181;182;186m&[0m[38;2;15;15;16m:[0m[38;2;19;19;19m:[0m[38;2;103;103;103m;[0m[38;2;187;187;187m;[0m[38;2;251;251;251m,[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m.[0m[38;2;255;255;255m.[0m[38;2;255;255;255m.[0m[38;2;255;255;255m,[0m[38;2;112;112;112ms[0m[38;2;0;0;0m.[0m[38;2;70;79;94m3[0m[38;2;128;145;171m9[0m[38;2;127;143;168m#[0m[38;2;127;143;168m#[0m[38;2;127;143;168m#[0m[38;2;127;143;168m#[0m[38;2;127;143;168m#[0m[38;2;127;143;168m#[0m[38;2;127;143;168m#[0m[38;2;127;143;168m#[0m[38;2;127;143;168m#[0m");
    $display("[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;235;235;235m:[0m[38;2;61;61;61mr[0m[38;2;0;0;0m.[0m[38;2;0;0;0m [0m[38;2;73;71;75m5[0m[38;2;242;226;217m@[0m[38;2;255;239;227m@[0m[38;2;255;238;227m@[0m[38;2;255;239;227m@[0m[38;2;255;242;231m@[0m[38;2;255;243;232m@[0m[38;2;221;206;198m@[0m[38;2;187;173;167mB[0m[38;2;170;158;152m9[0m[38;2;141;133;129m#[0m[38;2;90;86;86mh[0m[38;2;19;20;23m;[0m[38;2;0;0;0m [0m[38;2;39;37;38ms[0m[38;2;185;173;166mB[0m[38;2;255;238;226m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;255;237;226m@[0m[38;2;255;241;230m@[0m[38;2;255;237;226m@[0m[38;2;255;237;226m@[0m[38;2;255;240;229m@[0m[38;2;255;243;232m@[0m[38;2;254;237;226m@[0m[38;2;223;209;200m@[0m[38;2;158;150;145m9[0m[38;2;81;76;74m3[0m[38;2;50;39;39ms[0m[38;2;48;35;36ms[0m[38;2;18;17;19m:[0m[38;2;163;153;148m9[0m[38;2;255;238;227m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;250;228;217m@[0m[38;2;249;225;215m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;255;240;229m@[0m[38;2;160;144;137m9[0m[38;2;2;1;1m.[0m[38;2;78;78;81m3[0m[38;2;229;232;237m@[0m[38;2;237;240;245m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;240;243;248m@[0m[38;2;142;143;149m#[0m[38;2;0;0;0m.[0m[38;2;102;102;102ms[0m[38;2;255;255;255m,[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m.[0m[38;2;196;196;196m;[0m[38;2;110;110;110m;[0m[38;2;76;76;75m;[0m[38;2;82;82;82m:[0m[38;2;117;117;117m:[0m[38;2;96;96;95mr[0m[38;2;3;3;2m.[0m[38;2;46;51;59mA[0m[38;2;127;143;169m9[0m[38;2;129;145;170m9[0m[38;2;127;143;168m#[0m[38;2;127;143;168m#[0m[38;2;127;143;168m#[0m[38;2;127;143;168m#[0m[38;2;127;143;168m#[0m[38;2;127;143;168m#[0m[38;2;127;143;168m#[0m[38;2;127;143;168m#[0m");
    $display("[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m.[0m[38;2;119;119;119ms[0m[38;2;0;0;0m.[0m[38;2;0;0;0m [0m[38;2;62;60;62m2[0m[38;2;238;222;213m@[0m[38;2;255;238;226m@[0m[38;2;254;237;225m@[0m[38;2;185;171;164mB[0m[38;2;86;81;79m3[0m[38;2;70;66;65m5[0m[38;2;17;16;17m:[0m[38;2;23;22;23m;[0m[38;2;111;103;100mH[0m[38;2;118;110;106mG[0m[38;2;100;94;91mM[0m[38;2;84;79;77m3[0m[38;2;66;62;61m2[0m[38;2;72;68;66m5[0m[38;2;178;166;161mB[0m[38;2;254;237;226m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;255;238;227m@[0m[38;2;255;241;230m@[0m[38;2;243;226;216m@[0m[38;2;199;188;180m&[0m[38;2;137;132;126mS[0m[38;2;82;77;75m3[0m[38;2;55;42;43mX[0m[38;2;82;51;52m2[0m[38;2;152;98;98mG[0m[38;2;225;154;151mB[0m[38;2;171;122;119m#[0m[38;2;2;2;3m.[0m[38;2;129;122;119mS[0m[38;2;255;238;227m@[0m[38;2;254;236;225m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;254;236;225m@[0m[38;2;254;237;226m@[0m[38;2;255;238;227m@[0m[38;2;255;243;232m@[0m[38;2;253;234;223m@[0m[38;2;85;77;74m3[0m[38;2;0;0;0m [0m[38;2;133;134;138m#[0m[38;2;240;242;248m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;237;240;245m@[0m[38;2;231;234;239m@[0m[38;2;82;82;85mh[0m[38;2;0;0;0m.[0m[38;2;123;123;123ms[0m[38;2;242;242;242m,[0m[38;2;234;234;234m,[0m[38;2;221;221;220m:[0m[38;2;224;224;224m:[0m[38;2;252;252;252m,[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;247;247;247m,[0m[38;2;130;130;130mr[0m[38;2;11;11;11m:[0m[38;2;38;38;41mX[0m[38;2;117;116;124mS[0m[38;2;135;135;139m#[0m[38;2;97;97;99mH[0m[38;2;39;39;41ms[0m[38;2;0;0;0m [0m[38;2;9;10;13m,[0m[38;2;89;99;116mH[0m[38;2;127;143;168m#[0m[38;2;131;147;173m9[0m[38;2;128;144;169m9[0m[38;2;127;143;168m#[0m[38;2;127;143;168m#[0m[38;2;127;143;168m#[0m[38;2;127;143;168m#[0m[38;2;127;143;168m#[0m[38;2;127;143;168m#[0m");
    $display("[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;192;192;192mr[0m[38;2;18;18;18m;[0m[38;2;0;0;0m [0m[38;2;45;44;46mX[0m[38;2;228;211;202m@[0m[38;2;255;238;227m@[0m[38;2;253;236;225m@[0m[38;2;246;228;218m@[0m[38;2;194;182;174m&[0m[38;2;119;112;109mG[0m[38;2;33;31;31mr[0m[38;2;16;16;16m:[0m[38;2;174;163;156mB[0m[38;2;255;250;238m@[0m[38;2;255;248;236m@[0m[38;2;255;240;229m@[0m[38;2;253;235;225m@[0m[38;2;255;237;226m@[0m[38;2;255;238;227m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;254;238;226m@[0m[38;2;212;198;190m&[0m[38;2;107;100;97mH[0m[38;2;66;57;57m2[0m[38;2;71;47;48mA[0m[38;2;103;62;62m3[0m[38;2;160;95;95mG[0m[38;2;217;144;141mB[0m[38;2;250;177;173m&[0m[38;2;255;186;183m@[0m[38;2;227;162;159m&[0m[38;2;65;49;50mA[0m[38;2;53;52;53mA[0m[38;2;214;198;190m@[0m[38;2;255;238;227m@[0m[38;2;253;235;224m@[0m[38;2;254;236;225m@[0m[38;2;255;238;227m@[0m[38;2;255;241;230m@[0m[38;2;255;243;232m@[0m[38;2;255;239;228m@[0m[38;2;235;219;209m@[0m[38;2;191;178;170m&[0m[38;2;111;101;97mH[0m[38;2;11;9;9m,[0m[38;2;25;25;27mi[0m[38;2;194;196;201m&[0m[38;2;240;243;248m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;240;243;248m@[0m[38;2;196;198;204m&[0m[38;2;22;22;24m;[0m[38;2;0;0;0m [0m[38;2;16;16;15m,[0m[38;2;41;41;41m;[0m[38;2;32;33;34m:[0m[38;2;22;24;26m:[0m[38;2;20;20;21m:[0m[38;2;76;76;76mi[0m[38;2;201;201;201mi[0m[38;2;235;235;235m:[0m[38;2;101;101;101mr[0m[38;2;0;0;0m,[0m[38;2;68;67;73m5[0m[38;2;175;172;186mB[0m[38;2;194;190;206m&[0m[38;2;209;208;219m@[0m[38;2;255;255;255m@[0m[38;2;237;237;238m@[0m[38;2;153;153;154m9[0m[38;2;67;67;68m5[0m[38;2;15;16;17m:[0m[38;2;32;35;42mr[0m[38;2;87;96;115mM[0m[38;2;126;141;167m#[0m[38;2;130;146;172m9[0m[38;2;127;143;168m#[0m[38;2;127;143;168m#[0m[38;2;127;143;168m#[0m[38;2;127;143;168m#[0m[38;2;127;143;168m#[0m");
    $display("[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;243;243;243m:[0m[38;2;76;76;76mr[0m[38;2;0;0;0m [0m[38;2;26;26;26mi[0m[38;2;202;189;181m&[0m[38;2;255;239;228m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;238;221;211m@[0m[38;2;232;216;207m@[0m[38;2;198;186;180m&[0m[38;2;89;84;83mh[0m[38;2;22;22;23m;[0m[38;2;105;98;96mM[0m[38;2;197;184;176m&[0m[38;2;243;226;215m@[0m[38;2;255;240;229m@[0m[38;2;255;244;233m@[0m[38;2;255;241;230m@[0m[38;2;255;238;227m@[0m[38;2;255;236;225m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;255;239;228m@[0m[38;2;184;173;168mB[0m[38;2;30;31;32mr[0m[38;2;38;22;23mi[0m[38;2;132;77;78mM[0m[38;2;195;114;114m#[0m[38;2;239;161;158m&[0m[38;2;254;183;180m@[0m[38;2;251;181;178m@[0m[38;2;250;185;180m@[0m[38;2;195;162;156mB[0m[38;2;172;161;155mB[0m[38;2;238;222;212m@[0m[38;2;255;245;233m@[0m[38;2;255;243;232m@[0m[38;2;255;241;230m@[0m[38;2;249;231;221m@[0m[38;2;225;210;201m@[0m[38;2;189;177;170m&[0m[38;2;136;130;127mS[0m[38;2;81;78;78m3[0m[38;2;35;33;33mr[0m[38;2;5;5;5m.[0m[38;2;0;1;1m.[0m[38;2;0;0;0m [0m[38;2;68;68;72m5[0m[38;2;227;229;235m@[0m[38;2;237;240;245m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;241;244;249m@[0m[38;2;155;156;162m9[0m[38;2;8;8;9m,[0m[38;2;0;0;0m [0m[38;2;17;22;29m;[0m[38;2;29;44;59mX[0m[38;2;31;46;62mX[0m[38;2;38;55;73mA[0m[38;2;31;41;55ms[0m[38;2;5;6;9m:[0m[38;2;22;21;21m:[0m[38;2;47;47;46m;[0m[38;2;3;3;3m,[0m[38;2;82;82;89mh[0m[38;2;183;180;195m&[0m[38;2;191;186;203m&[0m[38;2;186;182;198m&[0m[38;2;196;194;207m&[0m[38;2;248;248;249m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;252;252;252m@[0m[38;2;204;204;206m@[0m[38;2;130;130;132mS[0m[38;2;43;43;44ms[0m[38;2;38;43;51ms[0m[38;2;102;115;137mG[0m[38;2;131;147;173m9[0m[38;2;129;145;170m9[0m[38;2;127;143;168m#[0m[38;2;127;143;168m#[0m[38;2;127;143;168m#[0m");
    $display("[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m.[0m[38;2;173;173;173mr[0m[38;2;12;12;12m:[0m[38;2;12;13;15m:[0m[38;2;191;180;175m&[0m[38;2;255;243;232m@[0m[38;2;255;237;225m@[0m[38;2;253;234;223m@[0m[38;2;195;182;175m&[0m[38;2;118;112;110mG[0m[38;2;70;67;67m5[0m[38;2;54;48;48mX[0m[38;2;17;15;16m:[0m[38;2;0;0;0m [0m[38;2;6;7;7m,[0m[38;2;36;35;35mr[0m[38;2;75;73;71m5[0m[38;2;135;127;123mS[0m[38;2;192;179;171m&[0m[38;2;231;214;205m@[0m[38;2;248;231;221m@[0m[38;2;255;240;229m@[0m[38;2;255;243;231m@[0m[38;2;255;244;232m@[0m[38;2;255;243;231m@[0m[38;2;255;242;230m@[0m[38;2;255;241;230m@[0m[38;2;255;240;229m@[0m[38;2;255;240;229m@[0m[38;2;255;239;228m@[0m[38;2;255;238;227m@[0m[38;2;255;238;227m@[0m[38;2;255;241;229m@[0m[38;2;236;219;209m@[0m[38;2;170;159;152m9[0m[38;2;121;115;111mG[0m[38;2;155;139;134m#[0m[38;2;241;209;199m@[0m[38;2;255;225;216m@[0m[38;2;255;229;219m@[0m[38;2;255;234;223m@[0m[38;2;253;235;224m@[0m[38;2;244;227;217m@[0m[38;2;215;201;192m@[0m[38;2;178;167;161mB[0m[38;2;137;130;125mS[0m[38;2;92;88;86mh[0m[38;2;57;55;55mA[0m[38;2;38;36;37mr[0m[38;2;44;34;34mr[0m[38;2;80;59;56m2[0m[38;2;103;74;69m3[0m[38;2;12;9;9m,[0m[38;2;7;8;8m,[0m[38;2;2;2;2m.[0m[38;2;14;14;15m:[0m[38;2;142;143;148m#[0m[38;2;236;239;244m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;236;239;244m@[0m[38;2;230;233;238m@[0m[38;2;86;86;90mh[0m[38;2;0;0;0m [0m[38;2;5;5;7m.[0m[38;2;33;46;62mX[0m[38;2;38;58;78mA[0m[38;2;53;71;89m5[0m[38;2;76;100;119mM[0m[38;2;77;101;120mM[0m[38;2;71;92;108mh[0m[38;2;37;48;57mX[0m[38;2;2;3;4m,[0m[38;2;3;2;2m.[0m[38;2;71;71;75m5[0m[38;2;154;151;164m9[0m[38;2;191;187;203m&[0m[38;2;189;185;202m&[0m[38;2;210;210;219m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;231;231;232m@[0m[38;2;115;115;115mG[0m[38;2;23;24;27mi[0m[38;2;61;68;81m5[0m[38;2;118;134;157m#[0m[38;2;131;147;173m9[0m[38;2;127;143;169m9[0m[38;2;127;143;168m#[0m");
    $display("[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;240;240;240m:[0m[38;2;63;63;63mr[0m[38;2;0;0;0m.[0m[38;2;113;107;105mH[0m[38;2;230;215;206m@[0m[38;2;250;232;222m@[0m[38;2;255;241;230m@[0m[38;2;255;247;235m@[0m[38;2;255;243;231m@[0m[38;2;241;224;214m@[0m[38;2;218;188;178m&[0m[38;2;202;154;142mB[0m[38;2;187;140;128m9[0m[38;2;181;133;122m#[0m[38;2;156;113;103mS[0m[38;2;95;69;63m3[0m[38;2;42;31;29mr[0m[38;2;21;16;17m:[0m[38;2;31;28;28mi[0m[38;2;54;51;50mA[0m[38;2;83;77;74m3[0m[38;2;112;104;99mH[0m[38;2;140;129;122mS[0m[38;2;163;151;145m9[0m[38;2;189;175;167mB[0m[38;2;198;183;176m&[0m[38;2;205;191;183m&[0m[38;2;207;193;185m&[0m[38;2;214;199;191m@[0m[38;2;227;211;201m@[0m[38;2;228;212;202m@[0m[38;2;225;209;199m@[0m[38;2;222;206;197m@[0m[38;2;216;201;193m@[0m[38;2;207;192;184m&[0m[38;2;194;181;172m&[0m[38;2;171;161;155mB[0m[38;2;148;139;133m#[0m[38;2;121;114;110mG[0m[38;2;89;84;80mh[0m[38;2;56;52;51mA[0m[38;2;38;35;35mr[0m[38;2;39;34;34mr[0m[38;2;52;40;39ms[0m[38;2;81;60;56m2[0m[38;2;122;91;86mM[0m[38;2;173;125;115m#[0m[38;2;210;156;142mB[0m[38;2;238;175;159m&[0m[38;2;255;190;171m@[0m[38;2;254;185;168m@[0m[38;2;101;77;73mh[0m[38;2;4;5;5m.[0m[38;2;13;13;13m:[0m[38;2;152;154;158m9[0m[38;2;240;243;248m@[0m[38;2;236;239;244m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;240;243;248m@[0m[38;2;181;183;187m&[0m[38;2;19;19;20m;[0m[38;2;0;0;0m [0m[38;2;21;28;38mi[0m[38;2;38;56;76mA[0m[38;2;41;59;77m2[0m[38;2;69;90;108mh[0m[38;2;79;105;125mH[0m[38;2;78;105;124mH[0m[38;2;79;106;125mH[0m[38;2;80;107;126mH[0m[38;2;66;85;101mh[0m[38;2;26;34;40mr[0m[38;2;0;0;0m [0m[38;2;11;11;11m,[0m[38;2;85;84;90mh[0m[38;2;140;138;149m#[0m[38;2;86;86;90mh[0m[38;2;186;187;190m&[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;186;186;187m&[0m[38;2;46;46;47mX[0m[38;2;21;25;30mi[0m[38;2;91;101;119mH[0m[38;2;129;145;171m9[0m[38;2;129;145;170m9[0m");
    $display("[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m.[0m[38;2;253;253;253m,[0m[38;2;238;238;238m,[0m[38;2;213;213;213m:[0m[38;2;161;161;161mr[0m[38;2;45;45;45m;[0m[38;2;0;0;0m.[0m[38;2;30;29;29mi[0m[38;2;65;62;61m2[0m[38;2;98;92;90mM[0m[38;2;132;123;119mS[0m[38;2;170;158;152m9[0m[38;2;204;190;183m&[0m[38;2;233;217;208m@[0m[38;2;253;231;220m@[0m[38;2;255;233;220m@[0m[38;2;255;225;210m@[0m[38;2;255;209;193m@[0m[38;2;255;197;180m@[0m[38;2;247;182;165m&[0m[38;2;207;148;136mB[0m[38;2;70;51;50mA[0m[38;2;0;0;0m [0m[38;2;0;0;3m.[0m[38;2;32;37;48ms[0m[38;2;24;27;32mi[0m[38;2;1;1;2m.[0m[38;2;0;0;0m [0m[38;2;0;0;0m [0m[38;2;1;1;1m.[0m[38;2;8;8;9m,[0m[38;2;25;25;26m;[0m[38;2;47;46;46ms[0m[38;2;55;53;52ms[0m[38;2;51;49;49mr[0m[38;2;47;46;46mi[0m[38;2;36;36;36mi[0m[38;2;20;19;20m:[0m[38;2;5;5;5m.[0m[38;2;0;0;0m [0m[38;2;0;0;0m [0m[38;2;0;0;0m [0m[38;2;0;0;0m [0m[38;2;0;0;0m [0m[38;2;36;29;28mr[0m[38;2;206;151;139mB[0m[38;2;247;182;165m&[0m[38;2;255;189;171m@[0m[38;2;255;192;173m@[0m[38;2;255;192;173m@[0m[38;2;255;189;171m@[0m[38;2;255;188;170m@[0m[38;2;255;190;172m@[0m[38;2;240;178;164m&[0m[38;2;85;66;63m5[0m[38;2;0;0;0m [0m[38;2;110;110;114mG[0m[38;2;237;239;245m@[0m[38;2;236;240;245m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;236;239;244m@[0m[38;2;235;238;243m@[0m[38;2;96;97;101mM[0m[38;2;0;0;0m [0m[38;2;10;13;18m:[0m[38;2;35;52;70mA[0m[38;2;37;57;76mA[0m[38;2;55;75;94m5[0m[38;2;78;104;123mH[0m[38;2;78;104;123mH[0m[38;2;78;104;123mH[0m[38;2;78;104;123mH[0m[38;2;78;104;123mH[0m[38;2;80;107;126mH[0m[38;2;75;99;117mM[0m[38;2;36;46;57mX[0m[38;2;6;8;12m,[0m[38;2;0;0;0m [0m[38;2;14;14;14m:[0m[38;2;0;0;0m [0m[38;2;40;40;43ms[0m[38;2;219;220;223m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;227;227;228m@[0m[38;2;91;91;92mh[0m[38;2;7;7;8m,[0m[38;2;61;68;80m5[0m[38;2;120;135;160m#[0m");
    $display("[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;247;247;247m,[0m[38;2;139;139;139mi[0m[38;2;60;60;60m:[0m[38;2;34;34;34m:[0m[38;2;26;26;27m;[0m[38;2;69;69;70ms[0m[38;2;58;58;58mr[0m[38;2;0;0;0m [0m[38;2;0;0;0m [0m[38;2;31;32;32m;[0m[38;2;41;42;43mr[0m[38;2;63;61;62m2[0m[38;2;63;60;60m2[0m[38;2;44;43;44ms[0m[38;2;42;41;42ms[0m[38;2;56;55;55mA[0m[38;2;88;84;82mh[0m[38;2;158;150;145m9[0m[38;2;242;227;217m@[0m[38;2;253;233;222m@[0m[38;2;255;226;213m@[0m[38;2;196;163;154mB[0m[38;2;22;18;18m;[0m[38;2;0;0;0m [0m[38;2;51;59;70m2[0m[38;2;132;146;171m9[0m[38;2;194;199;209m@[0m[38;2;184;185;189m&[0m[38;2;136;137;141m#[0m[38;2;103;103;107mH[0m[38;2;72;72;75m5[0m[38;2;42;42;44ms[0m[38;2;21;21;22m;[0m[38;2;33;33;33m;[0m[38;2;97;97;97mr[0m[38;2;130;130;131ms[0m[38;2;88;88;89mX[0m[38;2;45;45;44mi[0m[38;2;15;15;14m,[0m[38;2;6;7;7m,[0m[38;2;12;13;19m:[0m[38;2;24;26;38mi[0m[38;2;32;33;51ms[0m[38;2;9;10;14m,[0m[38;2;0;0;0m [0m[38;2;63;47;46mA[0m[38;2;245;179;164m&[0m[38;2;255;191;173m@[0m[38;2;254;186;169m@[0m[38;2;254;186;168m@[0m[38;2;254;186;169m@[0m[38;2;254;186;169m@[0m[38;2;255;191;173m@[0m[38;2;223;166;152m&[0m[38;2;80;60;56m2[0m[38;2;0;0;0m [0m[38;2;84;85;88mh[0m[38;2;225;228;232m@[0m[38;2;238;241;246m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;240;243;248m@[0m[38;2;186;188;194m&[0m[38;2;24;24;25m;[0m[38;2;0;0;0m [0m[38;2;27;37;49ms[0m[38;2;38;58;78mA[0m[38;2;44;62;80m2[0m[38;2;72;95;114mM[0m[38;2;79;105;124mH[0m[38;2;78;104;123mH[0m[38;2;78;104;123mH[0m[38;2;78;104;123mH[0m[38;2;78;104;123mH[0m[38;2;78;104;123mH[0m[38;2;79;105;124mH[0m[38;2;62;83;101m3[0m[38;2;36;52;69mA[0m[38;2;22;30;39mi[0m[38;2;4;5;8m.[0m[38;2;0;0;0m [0m[38;2;3;3;3m.[0m[38;2;165;166;170mB[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;251;251;252m@[0m[38;2;146;146;148m9[0m[38;2;15;14;15m:[0m[38;2;31;35;42mr[0m");
    $display("[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;182;182;182mr[0m[38;2;8;8;8m:[0m[38;2;0;0;0m [0m[38;2;53;53;56mA[0m[38;2;147;145;157m9[0m[38;2;167;164;178mB[0m[38;2;146;144;156m9[0m[38;2;120;120;130mS[0m[38;2;50;50;54mX[0m[38;2;0;0;0m [0m[38;2;50;48;48mX[0m[38;2;221;205;197m@[0m[38;2;253;236;225m@[0m[38;2;234;218;209m@[0m[38;2;211;196;188m&[0m[38;2;178;166;160mB[0m[38;2;146;137;132m#[0m[38;2;163;153;148m9[0m[38;2;240;224;214m@[0m[38;2;255;238;227m@[0m[38;2;255;241;230m@[0m[38;2;154;146;142m9[0m[38;2;9;8;8m,[0m[38;2;29;33;40mr[0m[38;2;118;131;153m#[0m[38;2;198;204;215m@[0m[38;2;238;240;245m@[0m[38;2;241;244;249m@[0m[38;2;243;246;251m@[0m[38;2;242;245;251m@[0m[38;2;238;240;246m@[0m[38;2;225;228;233m@[0m[38;2;197;199;204m&[0m[38;2;115;116;120mG[0m[38;2;2;2;3m.[0m[38;2;0;0;0m [0m[38;2;0;0;0m [0m[38;2;12;13;22m:[0m[38;2;40;40;69mX[0m[38;2;61;59;101m5[0m[38;2;70;67;115mh[0m[38;2;73;69;121mh[0m[38;2;75;71;124mh[0m[38;2;56;57;96m5[0m[38;2;16;17;26m;[0m[38;2;16;11;10m:[0m[38;2;124;90;86mM[0m[38;2;237;174;159m&[0m[38;2;255;192;173m@[0m[38;2;255;187;169m@[0m[38;2;255;187;169m@[0m[38;2;255;191;173m@[0m[38;2;199;145;133m9[0m[38;2;48;37;36ms[0m[38;2;0;0;0m [0m[38;2;78;78;81m3[0m[38;2;219;222;227m@[0m[38;2;239;242;247m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;236;240;245m@[0m[38;2;232;235;240m@[0m[38;2;92;92;95mM[0m[38;2;0;0;0m [0m[38;2;0;0;0m [0m[38;2;27;35;45mr[0m[38;2;40;60;80m2[0m[38;2;64;85;104mh[0m[38;2;81;107;126mH[0m[38;2;78;104;123mH[0m[38;2;78;104;123mH[0m[38;2;78;104;123mH[0m[38;2;78;104;123mH[0m[38;2;78;104;123mH[0m[38;2;78;104;123mH[0m[38;2;79;105;124mH[0m[38;2;74;96;114mM[0m[38;2;44;63;81m2[0m[38;2;38;57;77mA[0m[38;2;16;20;28m;[0m[38;2;0;0;0m [0m[38;2;12;12;14m:[0m[38;2;184;185;189m&[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;176;176;178mB[0m[38;2;23;23;23m;[0m");
    $display("[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;191;191;191mr[0m[38;2;14;14;14m:[0m[38;2;1;1;2m.[0m[38;2;160;160;166mB[0m[38;2;191;191;197m&[0m[38;2;79;78;85m3[0m[38;2;123;121;131mS[0m[38;2;172;170;183mB[0m[38;2;70;70;75m5[0m[38;2;1;1;1m.[0m[38;2;135;127;124mS[0m[38;2;255;238;227m@[0m[38;2;255;237;225m@[0m[38;2;255;238;226m@[0m[38;2;255;240;228m@[0m[38;2;255;242;230m@[0m[38;2;255;243;232m@[0m[38;2;255;242;230m@[0m[38;2;254;236;225m@[0m[38;2;255;241;230m@[0m[38;2;190;178;172m&[0m[38;2;24;24;24m;[0m[38;2;15;18;22m;[0m[38;2;113;123;141mS[0m[38;2;207;212;223m@[0m[38;2;242;245;249m@[0m[38;2;240;243;248m@[0m[38;2;239;242;247m@[0m[38;2;239;242;247m@[0m[38;2;238;241;246m@[0m[38;2;237;240;245m@[0m[38;2;237;240;245m@[0m[38;2;241;244;249m@[0m[38;2;236;238;244m@[0m[38;2;143;144;147m#[0m[38;2;45;45;47mX[0m[38;2;1;1;1m.[0m[38;2;13;14;22m:[0m[38;2;36;37;61mX[0m[38;2;55;54;92m5[0m[38;2;72;72;116mh[0m[38;2;86;87;131mH[0m[38;2;92;96;137mH[0m[38;2;99;104;145mG[0m[38;2;93;97;134mH[0m[38;2;46;50;65mA[0m[38;2;1;4;7m.[0m[38;2;54;39;37ms[0m[38;2;181;131;120m#[0m[38;2;253;185;168m@[0m[38;2;255;188;171m@[0m[38;2;159;118;111mS[0m[38;2;26;20;20m;[0m[38;2;0;0;0m [0m[38;2;83;84;87mh[0m[38;2;219;222;227m@[0m[38;2;239;243;248m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;241;244;250m@[0m[38;2;170;170;175mB[0m[38;2;15;15;15m:[0m[38;2;1;1;1m.[0m[38;2;2;2;2m.[0m[38;2;22;28;36mi[0m[38;2;28;38;51ms[0m[38;2;40;50;61mX[0m[38;2;66;86;102mh[0m[38;2;80;106;126mH[0m[38;2;79;106;125mH[0m[38;2;78;104;123mH[0m[38;2;78;104;123mH[0m[38;2;78;104;123mH[0m[38;2;78;104;123mH[0m[38;2;78;104;123mH[0m[38;2;79;104;123mH[0m[38;2;60;80;97m3[0m[38;2;37;52;70mA[0m[38;2;10;12;15m:[0m[38;2;0;0;0m [0m[38;2;100;101;104mH[0m[38;2;248;248;249m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;168;168;171mB[0m");
    $display("[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;197;197;197mr[0m[38;2;15;15;16m:[0m[38;2;38;38;40ms[0m[38;2;220;221;223m@[0m[38;2;247;248;248m@[0m[38;2;134;134;136m#[0m[38;2;20;20;21m;[0m[38;2;13;14;15m:[0m[38;2;3;3;4m.[0m[38;2;67;63;62m2[0m[38;2;242;225;215m@[0m[38;2;255;240;229m@[0m[38;2;253;236;225m@[0m[38;2;253;236;225m@[0m[38;2;253;236;225m@[0m[38;2;253;236;226m@[0m[38;2;253;237;226m@[0m[38;2;253;237;226m@[0m[38;2;255;241;230m@[0m[38;2;215;200;193m@[0m[38;2;47;45;45mX[0m[38;2;2;4;5m.[0m[38;2;87;95;109mM[0m[38;2;180;185;195m&[0m[38;2;206;209;213m@[0m[38;2;199;202;207m@[0m[38;2;197;199;205m&[0m[38;2;200;202;207m@[0m[38;2;206;209;213m@[0m[38;2;219;221;226m@[0m[38;2;233;236;241m@[0m[38;2;242;245;250m@[0m[38;2;239;242;247m@[0m[38;2;236;239;244m@[0m[38;2;245;248;253m@[0m[38;2;196;198;203m&[0m[38;2;33;33;35mr[0m[38;2;0;0;0m [0m[38;2;1;0;0m.[0m[38;2;0;0;0m [0m[38;2;12;14;18m:[0m[38;2;35;38;46ms[0m[38;2;60;64;83m5[0m[38;2;85;90;119mM[0m[38;2;99;106;144mG[0m[38;2;107;115;152mS[0m[38;2;85;91;120mM[0m[38;2;34;37;54ms[0m[38;2;14;13;16m:[0m[38;2;81;60;56m2[0m[38;2;99;75;70m3[0m[38;2;6;6;6m,[0m[38;2;0;0;0m [0m[38;2;92;93;96mM[0m[38;2;219;221;226m@[0m[38;2;237;240;246m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;239;242;247m@[0m[38;2;212;214;220m@[0m[38;2;54;53;55mA[0m[38;2;3;3;3m.[0m[38;2;6;6;6m.[0m[38;2;7;7;9m,[0m[38;2;29;40;53ms[0m[38;2;22;32;42mr[0m[38;2;9;12;16m:[0m[38;2;8;9;10m,[0m[38;2;33;42;50ms[0m[38;2;68;89;107mh[0m[38;2;80;107;127mH[0m[38;2;79;105;124mH[0m[38;2;78;104;123mH[0m[38;2;78;104;123mH[0m[38;2;78;104;123mH[0m[38;2;78;105;124mH[0m[38;2;76;98;117mM[0m[38;2;40;50;63mX[0m[38;2;1;1;2m.[0m[38;2;31;32;33mr[0m[38;2;216;216;218m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m");
    $display("[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m.[0m[38;2;131;131;131ms[0m[38;2;0;0;0m.[0m[38;2;103;104;108mH[0m[38;2;251;252;253m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;200;200;201m&[0m[38;2;69;70;72m5[0m[38;2;4;4;5m.[0m[38;2;33;30;30mr[0m[38;2;163;151;145m9[0m[38;2;242;223;213m@[0m[38;2;255;237;225m@[0m[38;2;255;234;222m@[0m[38;2;255;232;220m@[0m[38;2;255;229;216m@[0m[38;2;255;225;211m@[0m[38;2;255;220;205m@[0m[38;2;235;193;180m@[0m[38;2;73;64;63m2[0m[38;2;0;0;0m [0m[38;2;14;15;17m:[0m[38;2;23;24;27mi[0m[38;2;24;24;25m;[0m[38;2;22;22;25m;[0m[38;2;35;37;42ms[0m[38;2;35;36;42ms[0m[38;2;34;35;40mr[0m[38;2;34;35;38mr[0m[38;2;39;39;42ms[0m[38;2;58;58;61m2[0m[38;2;112;112;114mG[0m[38;2;203;205;209m@[0m[38;2;238;241;246m@[0m[38;2;237;241;246m@[0m[38;2;223;225;232m@[0m[38;2;66;66;70m5[0m[38;2;0;0;0m [0m[38;2;24;30;39mr[0m[38;2;17;22;31m;[0m[38;2;3;3;5m.[0m[38;2;1;0;0m.[0m[38;2;4;4;3m.[0m[38;2;10;10;13m,[0m[38;2;19;20;29m;[0m[38;2;37;39;51ms[0m[38;2;55;58;75m2[0m[38;2;56;59;80m2[0m[38;2;35;37;49ms[0m[38;2;7;10;11m,[0m[38;2;0;0;0m [0m[38;2;0;0;0m [0m[38;2;64;64;66m2[0m[38;2;199;200;209m@[0m[38;2;224;226;232m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;238;241;245m@[0m[38;2;226;230;237m@[0m[38;2;95;98;107mM[0m[38;2;0;0;0m [0m[38;2;16;16;18m:[0m[38;2;3;2;2m.[0m[38;2;17;20;26m;[0m[38;2;44;60;78m2[0m[38;2;39;58;78mA[0m[38;2;37;56;74mA[0m[38;2;30;43;58ms[0m[38;2;11;14;19m:[0m[38;2;9;11;14m,[0m[38;2;44;58;71mA[0m[38;2;76;100;119mM[0m[38;2;80;106;125mH[0m[38;2;79;106;125mH[0m[38;2;79;106;125mH[0m[38;2;79;106;125mH[0m[38;2;79;104;123mH[0m[38;2;32;39;46ms[0m[38;2;0;0;0m [0m[38;2;116;116;120mG[0m[38;2;253;253;253m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m");
    $display("[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;240;240;240m:[0m[38;2;63;63;63mr[0m[38;2;7;7;8m,[0m[38;2;174;174;177mB[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;251;251;252m@[0m[38;2;193;194;195m&[0m[38;2;100;101;102mM[0m[38;2;23;24;25m;[0m[38;2;44;37;36ms[0m[38;2;127;96;90mH[0m[38;2;181;137;125m9[0m[38;2;183;138;125m9[0m[38;2;167;121;111mS[0m[38;2;146;103;94mG[0m[38;2;124;88;80mM[0m[38;2;57;42;39mX[0m[38;2;0;0;0m [0m[38;2;14;14;15m:[0m[38;2;29;29;32mi[0m[38;2;1;1;1m.[0m[38;2;0;0;0m [0m[38;2;11;11;13m,[0m[38;2;94;104;122mH[0m[38;2;121;136;160m#[0m[38;2;117;131;154m#[0m[38;2;111;125;148mS[0m[38;2;96;109;132mG[0m[38;2;75;86;104mh[0m[38;2;43;50;62mA[0m[38;2;77;80;88m3[0m[38;2;210;213;219m@[0m[38;2;240;243;248m@[0m[38;2;218;220;227m@[0m[38;2;59;59;62m2[0m[38;2;0;0;0m [0m[38;2;32;44;59mX[0m[38;2;31;43;59ms[0m[38;2;20;25;34mi[0m[38;2;17;22;30m;[0m[38;2;3;3;3m.[0m[38;2;10;11;15m:[0m[38;2;29;33;54ms[0m[38;2;34;36;62ms[0m[38;2;21;23;39mi[0m[38;2;16;18;30m;[0m[38;2;24;26;42mi[0m[38;2;15;15;18m:[0m[38;2;0;0;0m [0m[38;2;61;60;62m2[0m[38;2;169;172;181mB[0m[38;2;195;199;210m@[0m[38;2;234;237;242m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;237;240;245m@[0m[38;2;228;231;238m@[0m[38;2;135;140;155m#[0m[38;2;12;13;16m:[0m[38;2;13;17;24m:[0m[38;2;12;13;17m:[0m[38;2;1;1;1m.[0m[38;2;43;54;66mA[0m[38;2;74;96;114mM[0m[38;2;53;71;89m5[0m[38;2;38;56;75mA[0m[38;2;39;58;78mA[0m[38;2;38;55;73mA[0m[38;2;21;27;36mi[0m[38;2;4;3;3m.[0m[38;2;20;25;30mi[0m[38;2;48;63;79m2[0m[38;2;60;81;100m3[0m[38;2;65;87;106mh[0m[38;2;71;95;114mM[0m[38;2;65;82;98m3[0m[38;2;9;11;14m,[0m[38;2;28;27;28mi[0m[38;2;206;205;207m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m");
    $display("[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;195;195;195mr[0m[38;2;15;15;15m:[0m[38;2;48;47;50mX[0m[38;2;227;227;229m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;220;220;221m@[0m[38;2;139;140;142m#[0m[38;2;72;74;76m5[0m[38;2;55;55;57mA[0m[38;2;59;58;60m2[0m[38;2;70;71;74m5[0m[38;2;91;94;96mM[0m[38;2;108;111;114mH[0m[38;2;135;137;139m#[0m[38;2;168;169;170mB[0m[38;2;178;179;182m&[0m[38;2;53;54;57mA[0m[38;2;2;2;3m.[0m[38;2;21;21;24m;[0m[38;2;2;1;1m.[0m[38;2;75;82;98mh[0m[38;2;130;146;172m9[0m[38;2;126;142;168m#[0m[38;2;142;154;176m9[0m[38;2;169;178;195m&[0m[38;2;176;185;202m&[0m[38;2;190;197;211m&[0m[38;2;193;198;207m&[0m[38;2;212;214;221m@[0m[38;2;239;242;247m@[0m[38;2;194;196;200m&[0m[38;2;28;28;29mi[0m[38;2;4;6;8m,[0m[38;2;36;51;68mA[0m[38;2;21;28;36mi[0m[38;2;6;7;8m,[0m[38;2;20;23;29m;[0m[38;2;4;4;5m.[0m[38;2;13;15;17m:[0m[38;2;6;6;8m,[0m[38;2;32;32;53ms[0m[38;2;67;65;110m3[0m[38;2;77;74;128mM[0m[38;2;55;56;94m5[0m[38;2;6;7;10m,[0m[38;2;48;48;50mX[0m[38;2;185;186;194m&[0m[38;2;156;165;183mB[0m[38;2;200;203;212m@[0m[38;2;237;240;245m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;236;239;244m@[0m[38;2;230;233;239m@[0m[38;2;158;166;182mB[0m[38;2;40;45;52mX[0m[38;2;18;21;36mi[0m[38;2;32;39;60ms[0m[38;2;1;1;2m.[0m[38;2;21;25;30mi[0m[38;2;73;95;114mM[0m[38;2;80;107;126mH[0m[38;2;78;102;121mM[0m[38;2;58;78;97m3[0m[38;2;39;57;75mA[0m[38;2;38;57;76mA[0m[38;2;39;58;77mA[0m[38;2;30;41;55ms[0m[38;2;6;7;9m,[0m[38;2;4;5;6m.[0m[38;2;26;35;47mr[0m[38;2;38;57;76mA[0m[38;2;40;58;77mA[0m[38;2;20;25;32mi[0m[38;2;0;0;0m [0m[38;2;101;100;103mH[0m[38;2;252;252;253m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m");
    $display("[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m.[0m[38;2;136;136;136ms[0m[38;2;0;0;0m.[0m[38;2;109;108;112mH[0m[38;2;254;254;254m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;249;249;250m@[0m[38;2;250;250;250m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;211;211;213m@[0m[38;2;26;26;27mi[0m[38;2;30;30;32mi[0m[38;2;58;57;61mA[0m[38;2;0;0;0m [0m[38;2;66;71;89m3[0m[38;2;129;144;171m9[0m[38;2;125;140;165m#[0m[38;2;188;193;205m&[0m[38;2;240;242;246m@[0m[38;2;238;241;245m@[0m[38;2;241;243;248m@[0m[38;2;242;245;250m@[0m[38;2;238;241;245m@[0m[38;2;240;242;248m@[0m[38;2;132;133;137m#[0m[38;2;3;2;2m.[0m[38;2;16;20;27m;[0m[38;2;38;54;73mA[0m[38;2;15;19;24m;[0m[38;2;0;0;0m [0m[38;2;0;0;0m [0m[38;2;18;21;24m;[0m[38;2;69;88;104mh[0m[38;2;46;57;66mA[0m[38;2;6;6;6m,[0m[38;2;12;12;18m:[0m[38;2;47;50;80m2[0m[38;2;21;23;34mi[0m[38;2;8;7;7m,[0m[38;2;139;140;147m#[0m[38;2;162;172;192mB[0m[38;2;129;143;168m9[0m[38;2;198;202;211m@[0m[38;2;237;240;245m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;236;239;243m@[0m[38;2;179;185;200m&[0m[38;2;66;74;88m3[0m[38;2;24;26;41mi[0m[38;2;56;59;100m5[0m[38;2;15;17;26m;[0m[38;2;4;4;4m.[0m[38;2;57;72;84m5[0m[38;2;80;107;126mH[0m[38;2;78;104;123mH[0m[38;2;78;105;124mH[0m[38;2;79;104;123mH[0m[38;2;64;85;103mh[0m[38;2;41;59;77m2[0m[38;2;37;56;75mA[0m[38;2;39;59;78mA[0m[38;2;35;49;65mX[0m[38;2;13;16;21m:[0m[38;2;3;2;2m.[0m[38;2;23;31;41mr[0m[38;2;27;36;48mr[0m[38;2;0;0;0m [0m[38;2;22;22;24m;[0m[38;2;198;197;199m&[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m");
    $display("[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;242;242;242m:[0m[38;2;69;69;70mr[0m[38;2;7;7;8m,[0m[38;2;176;176;179mB[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;253;253;253m@[0m[38;2;113;112;115mG[0m[38;2;0;0;0m [0m[38;2;93;94;99mM[0m[38;2;76;77;82m3[0m[38;2;0;0;0m [0m[38;2;68;73;90m3[0m[38;2;126;142;169m#[0m[38;2;148;159;179mB[0m[38;2;223;225;232m@[0m[38;2;237;240;244m@[0m[38;2;237;240;245m@[0m[38;2;227;230;235m@[0m[38;2;216;219;224m@[0m[38;2;238;241;246m@[0m[38;2;216;219;224m@[0m[38;2;56;56;59mA[0m[38;2;2;2;3m.[0m[38;2;30;42;57ms[0m[38;2;37;55;75mA[0m[38;2;10;13;19m:[0m[38;2;0;0;0m [0m[38;2;8;10;12m,[0m[38;2;59;74;89m5[0m[38;2;80;107;126mH[0m[38;2;80;106;126mH[0m[38;2;62;80;95m3[0m[38;2;20;25;29mi[0m[38;2;3;4;4m.[0m[38;2;1;1;1m.[0m[38;2;56;56;58mA[0m[38;2;156;163;178mB[0m[38;2;78;88;104mh[0m[38;2;82;94;113mM[0m[38;2;189;197;210m&[0m[38;2;238;240;245m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;237;240;245m@[0m[38;2;204;209;219m@[0m[38;2;82;90;106mM[0m[38;2;12;14;19m:[0m[38;2;61;61;103m3[0m[38;2;37;39;64mX[0m[38;2;0;0;0m [0m[38;2;33;40;47ms[0m[38;2;78;102;121mM[0m[38;2;78;105;124mH[0m[38;2;78;104;123mH[0m[38;2;78;104;123mH[0m[38;2;78;104;123mH[0m[38;2;79;105;124mH[0m[38;2;70;91;109mh[0m[38;2;46;63;81m2[0m[38;2;37;56;75mA[0m[38;2;39;58;78mA[0m[38;2;38;55;74mA[0m[38;2;22;29;39mi[0m[38;2;2;2;2m.[0m[38;2;0;0;0m [0m[38;2;31;31;32mr[0m[38;2;174;174;176mB[0m[38;2;254;254;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;247;247;248m@[0m");
    $display("[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;199;199;199mr[0m[38;2;18;18;18m:[0m[38;2;48;48;51mX[0m[38;2;230;230;232m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;208;208;210m@[0m[38;2;27;27;29mi[0m[38;2;25;26;27mi[0m[38;2;146;145;155m9[0m[38;2;50;50;54mX[0m[38;2;1;2;2m.[0m[38;2;83;93;110mM[0m[38;2;140;153;176m9[0m[38;2;209;213;222m@[0m[38;2;238;240;245m@[0m[38;2;237;240;245m@[0m[38;2;223;226;231m@[0m[38;2;82;83;85mh[0m[38;2;30;30;32mi[0m[38;2;178;179;183m&[0m[38;2;163;164;169mB[0m[38;2;4;3;4m.[0m[38;2;9;12;16m:[0m[38;2;37;54;72mA[0m[38;2;33;48;64mX[0m[38;2;3;4;6m.[0m[38;2;12;14;16m:[0m[38;2;57;75;90m5[0m[38;2;79;106;126mH[0m[38;2;78;104;123mH[0m[38;2;78;104;123mH[0m[38;2;80;107;126mH[0m[38;2;76;101;120mM[0m[38;2;34;44;52ms[0m[38;2;1;1;1m.[0m[38;2;78;79;83m3[0m[38;2;70;73;82m3[0m[38;2;1;2;2m.[0m[38;2;36;41;49ms[0m[38;2;183;190;202m&[0m[38;2;238;241;246m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;236;239;244m@[0m[38;2;228;231;237m@[0m[38;2;130;138;154m#[0m[38;2;14;16;19m:[0m[38;2;23;24;37mi[0m[38;2;53;56;93m5[0m[38;2;7;7;10m,[0m[38;2;11;13;16m:[0m[38;2;67;87;103mh[0m[38;2;79;106;126mH[0m[38;2;78;104;123mH[0m[38;2;78;104;123mH[0m[38;2;78;104;123mH[0m[38;2;78;104;123mH[0m[38;2;78;104;123mH[0m[38;2;79;106;125mH[0m[38;2;74;96;115mM[0m[38;2;50;68;86m5[0m[38;2;38;58;78mA[0m[38;2;36;52;70mA[0m[38;2;17;22;30m;[0m[38;2;0;0;0m [0m[38;2;58;59;62m2[0m[38;2;206;207;209m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;242;242;243m@[0m[38;2;190;190;192m&[0m[38;2;109;109;111mH[0m[38;2;45;45;46mX[0m");
    $display("[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m.[0m[38;2;131;131;131ms[0m[38;2;0;0;0m.[0m[38;2;115;115;118mG[0m[38;2;253;253;254m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;252;252;252m@[0m[38;2;114;114;116mG[0m[38;2;0;0;0m [0m[38;2;93;93;100mM[0m[38;2;151;150;162m9[0m[38;2;16;16;16m:[0m[38;2;29;34;40mr[0m[38;2;130;142;162m#[0m[38;2;210;214;224m@[0m[38;2;242;245;248m@[0m[38;2;240;243;248m@[0m[38;2;242;245;250m@[0m[38;2;167;169;174mB[0m[38;2;8;8;9m,[0m[38;2;0;0;0m [0m[38;2;96;96;101mM[0m[38;2;98;99;104mM[0m[38;2;43;43;46ms[0m[38;2;7;7;8m,[0m[38;2;10;13;17m:[0m[38;2;9;10;13m,[0m[38;2;26;32;38mr[0m[38;2;67;88;105mh[0m[38;2;80;106;126mH[0m[38;2;78;104;123mH[0m[38;2;78;104;123mH[0m[38;2;78;104;123mH[0m[38;2;78;104;123mH[0m[38;2;81;107;127mH[0m[38;2;52;66;78m2[0m[38;2;5;5;5m.[0m[38;2;23;23;26m;[0m[38;2;4;4;5m.[0m[38;2;0;0;0m [0m[38;2;20;22;28m;[0m[38;2;176;181;193m&[0m[38;2;241;244;248m@[0m[38;2;236;239;244m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;238;241;245m@[0m[38;2;196;202;212m@[0m[38;2;67;75;89m3[0m[38;2;0;0;0m [0m[38;2;30;33;51ms[0m[38;2;25;27;42mr[0m[38;2;1;0;0m.[0m[38;2;46;57;69mA[0m[38;2;79;105;124mH[0m[38;2;78;104;123mH[0m[38;2;78;104;123mH[0m[38;2;78;104;123mH[0m[38;2;78;104;123mH[0m[38;2;78;104;123mH[0m[38;2;78;104;123mH[0m[38;2;78;105;124mH[0m[38;2;80;106;125mH[0m[38;2;72;93;111mM[0m[38;2;36;47;60mX[0m[38;2;5;7;12m,[0m[38;2;18;17;19m:[0m[38;2;125;125;127mS[0m[38;2;236;236;237m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;249;249;250m@[0m[38;2;202;202;203m@[0m[38;2;119;119;121mG[0m[38;2;46;47;49mX[0m[38;2;23;23;25m;[0m[38;2;54;53;58mA[0m[38;2;57;57;60mA[0m");
    $display("[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;238;238;238m:[0m[38;2;64;64;64mr[0m[38;2;10;11;11m:[0m[38;2;182;183;185m&[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;204;205;208m@[0m[38;2;29;29;31mi[0m[38;2;21;21;22m;[0m[38;2;158;156;168m9[0m[38;2;121;120;128mS[0m[38;2;23;26;30mi[0m[38;2;117;124;142mS[0m[38;2;197;201;213m@[0m[38;2;199;204;212m@[0m[38;2;167;171;179mB[0m[38;2;123;125;133mS[0m[38;2;88;89;93mh[0m[38;2;40;41;43ms[0m[38;2;18;18;21m;[0m[38;2;22;22;24m;[0m[38;2;79;78;83m3[0m[38;2;141;141;149m#[0m[38;2;193;192;203m&[0m[38;2;133;134;138m#[0m[38;2;27;27;28mi[0m[38;2;2;2;2m.[0m[38;2;41;52;62mA[0m[38;2;74;98;116mM[0m[38;2;78;104;123mH[0m[38;2;78;104;123mH[0m[38;2;78;104;123mH[0m[38;2;78;104;123mH[0m[38;2;78;104;123mH[0m[38;2;79;105;124mH[0m[38;2;72;94;112mM[0m[38;2;23;28;33mi[0m[38;2;0;0;0m [0m[38;2;12;14;18m:[0m[38;2;16;19;25m;[0m[38;2;12;13;14m:[0m[38;2;142;148;160m9[0m[38;2;214;218;227m@[0m[38;2;228;231;237m@[0m[38;2;234;237;242m@[0m[38;2;236;239;244m@[0m[38;2;232;235;240m@[0m[38;2;165;172;188mB[0m[38;2;53;57;66mA[0m[38;2;0;0;0m [0m[38;2;19;22;29m;[0m[38;2;2;3;3m.[0m[38;2;22;27;31mi[0m[38;2;75;97;115mM[0m[38;2;79;105;125mH[0m[38;2;78;104;123mH[0m[38;2;78;104;123mH[0m[38;2;78;104;123mH[0m[38;2;78;104;123mH[0m[38;2;78;104;123mH[0m[38;2;78;103;123mH[0m[38;2;72;94;112mM[0m[38;2;56;73;90m5[0m[38;2;29;35;43mr[0m[38;2;5;5;6m.[0m[38;2;54;53;55mA[0m[38;2;188;188;191m&[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;238;239;240m@[0m[38;2;169;169;171mB[0m[38;2;75;75;78m3[0m[38;2;17;17;19m:[0m[38;2;36;36;39mr[0m[38;2;102;101;108mH[0m[38;2;159;156;168mB[0m[38;2;189;185;200m&[0m[38;2;186;183;198m&[0m");

	$display("\033[31m \033[5m     //   / /     //   ) )     //   ) )     //   ) )     //   ) )\033[0m");
    $display("\033[31m \033[5m    //____       //___/ /     //___/ /     //   / /     //___/ /\033[0m");
    $display("\033[31m \033[5m   / ____       / ___ (      / ___ (      //   / /     / ___ (\033[0m");
    $display("\033[31m \033[5m  //           //   | |     //   | |     //   / /     //   | |\033[0m");
    $display("\033[31m \033[5m //____/ /    //    | |    //    | |    ((___/ /     //    | |\033[0m");
end endtask

task display_pass; begin
    $display("[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;254m.[0m[38;2;245;245;244m9[0m[38;2;187;187;188m&[0m[38;2;236;236;236m&[0m[38;2;255;255;254m;[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m;[0m[38;2;242;242;243m9[0m[38;2;175;174;175m&[0m[38;2;224;224;224mB[0m[38;2;255;255;255mX[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255ms[0m[38;2;214;214;215m&[0m[38;2;194;194;196m&[0m[38;2;255;255;255m3[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255mr[0m[38;2;217;217;217m9[0m[38;2;229;229;230m#[0m[38;2;255;255;255m,[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;251;251;251m5[0m[38;2;245;245;245m3[0m[38;2;255;254;254m,[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;253;253;253mS[0m[38;2;179;179;180m&[0m[38;2;219;219;220m&[0m[38;2;255;255;255mA[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255ms[0m[38;2;231;229;226m&[0m[38;2;220;215;208m@[0m[38;2;255;255;235mG[0m[38;2;251;238;212m3[0m[38;2;205;191;167mh[0m[38;2;154;142;121m3[0m[38;2;166;148;117mH[0m[38;2;202;177;128m9[0m[38;2;232;201;138m&[0m[38;2;252;219;150m&[0m[38;2;255;230;164m&[0m[38;2;255;237;184m9[0m[38;2;255;244;209mH[0m[38;2;255;250;232m2[0m[38;2;255;253;249m;[0m[38;2;255;255;255m.[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m");
    $display("[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m:[0m[38;2;250;250;250mA[0m[38;2;248;248;248mX[0m[38;2;255;255;255m,[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m:[0m[38;2;245;244;245m#[0m[38;2;182;181;183m&[0m[38;2;214;214;214mB[0m[38;2;255;255;255m5[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m.[0m[38;2;227;227;227m,[0m[38;2;177;177;176m:[0m[38;2;135;135;135m:[0m[38;2;120;119;121mi[0m[38;2;99;98;100m5[0m[38;2;72;72;73m3[0m[38;2;212;212;213mB[0m[38;2;255;255;255mi[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m.[0m[38;2;255;255;255m:[0m[38;2;255;255;255m:[0m[38;2;255;255;255m.[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255mr[0m[38;2;206;206;206m&[0m[38;2;209;209;210m&[0m[38;2;255;255;255m;[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;253;253;253mG[0m[38;2;184;184;186m&[0m[38;2;211;211;211m&[0m[38;2;255;255;255m5[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;252;245mi[0m[38;2;254;243;219mM[0m[38;2;254;238;204mG[0m[38;2;255;241;198m#[0m[38;2;248;225;177mB[0m[38;2;203;182;139m9[0m[38;2;144;128;94mH[0m[38;2;106;96;65m3[0m[38;2;127;119;71mH[0m[38;2;175;167;95m9[0m[38;2;147;139;80mS[0m[38;2;117;109;66mM[0m[38;2;101;93;58mh[0m[38;2;102;92;58mh[0m[38;2;121;106;70mM[0m[38;2;154;132;89mS[0m[38;2;190;165;111m9[0m[38;2;225;197;140mB[0m[38;2;250;224;172m9[0m[38;2;255;242;203mG[0m[38;2;255;251;228m5[0m[38;2;255;254;245mr[0m[38;2;255;255;253m,[0m[38;2;253;253;254ms[0m");
    $display("[38;2;225;225;225m#[0m[38;2;250;250;250m3[0m[38;2;254;254;254m:[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m,[0m[38;2;246;245;245mh[0m[38;2;243;243;242mh[0m[38;2;255;255;255m;[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m.[0m[38;2;251;251;251mG[0m[38;2;191;191;191m&[0m[38;2;211;211;212m&[0m[38;2;255;255;255m2[0m[38;2;249;249;249m.[0m[38;2;176;176;175m:[0m[38;2;88;88;88m;[0m[38;2;45;45;47mr[0m[38;2;42;42;46mX[0m[38;2;55;56;62m5[0m[38;2;63;63;70m5[0m[38;2;26;26;28mi[0m[38;2;3;3;3m.[0m[38;2;54;54;55m2[0m[38;2;234;234;234mS[0m[38;2;255;255;255m,[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;254;254;254mH[0m[38;2;178;178;180m&[0m[38;2;239;239;239m9[0m[38;2;255;255;255m.[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m,[0m[38;2;250;249;249mG[0m[38;2;185;185;186m&[0m[38;2;210;209;210m&[0m[38;2;255;255;255m5[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;253m2[0m[38;2;246;229;194mB[0m[38;2;250;218;150m@[0m[38;2;244;211;140m@[0m[38;2;144;124;83mG[0m[38;2;92;82;53m3[0m[38;2;119;111;65mM[0m[38;2;181;173;99m9[0m[38;2;233;224;126m&[0m[38;2;255;248;140m@[0m[38;2;255;251;142m@[0m[38;2;255;252;143m@[0m[38;2;255;249;141m@[0m[38;2;251;240;136m@[0m[38;2;231;221;125m&[0m[38;2;202;193;110mB[0m[38;2;164;157;90m#[0m[38;2;127;121;70mH[0m[38;2;101;94;56mh[0m[38;2;94;85;53m3[0m[38;2;119;103;68mM[0m[38;2;166;145;102mS[0m[38;2;220;196;147m#[0m[38;2;255;235;190m#[0m[38;2;255;240;210m&[0m");
    $display("[38;2;189;189;189mB[0m[38;2;178;178;179m&[0m[38;2;246;245;246mB[0m[38;2;253;253;253m,[0m[38;2;255;255;255m,[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;254;254;254m:[0m[38;2;238;238;239m9[0m[38;2;220;220;220mB[0m[38;2;255;255;254m2[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m2[0m[38;2;241;242;242mS[0m[38;2;196;195;194mH[0m[38;2;60;60;59m,[0m[38;2;20;21;23mi[0m[38;2;53;53;58m2[0m[38;2;78;78;85m3[0m[38;2;84;85;93mh[0m[38;2;83;83;91mh[0m[38;2;42;42;45ms[0m[38;2;41;42;45ms[0m[38;2;74;75;82m3[0m[38;2;16;17;19m;[0m[38;2;85;84;85m5[0m[38;2;183;183;183mX[0m[38;2;169;169;169m:[0m[38;2;169;169;169m:[0m[38;2;183;183;183m:[0m[38;2;234;234;234m,[0m[38;2;255;255;255m.[0m[38;2;255;255;255m.[0m[38;2;255;255;255m.[0m[38;2;255;255;255m.[0m[38;2;255;255;255m [0m[38;2;255;255;255mh[0m[38;2;232;232;232m9[0m[38;2;255;255;255mA[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m;[0m[38;2;249;249;249mA[0m[38;2;254;254;254mr[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255ms[0m[38;2;214;213;215m&[0m[38;2;209;209;209mB[0m[38;2;255;255;255m2[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255mr[0m[38;2;240;240;241m#[0m[38;2;204;199;194m&[0m[38;2;230;208;161m@[0m[38;2;254;222;148m@[0m[38;2;231;201;138m&[0m[38;2;19;17;14m:[0m[38;2;154;146;84mS[0m[38;2;255;255;145m@[0m[38;2;255;250;142m@[0m[38;2;255;245;139m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;244;138m@[0m[38;2;255;246;139m@[0m[38;2;255;248;141m@[0m[38;2;255;251;142m@[0m[38;2;255;251;142m@[0m[38;2;255;244;138m@[0m[38;2;232;223;126m&[0m[38;2;193;185;106mB[0m[38;2;137;131;75mG[0m[38;2;90;83;49m3[0m[38;2;93;81;53m3[0m[38;2;163;143;99mS[0m");
    $display("[38;2;255;255;255mr[0m[38;2;251;251;251mX[0m[38;2;253;253;253ms[0m[38;2;247;247;247mS[0m[38;2;208;208;209mB[0m[38;2;228;228;228m#[0m[38;2;251;251;251m5[0m[38;2;255;255;255m:[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m.[0m[38;2;255;255;255m.[0m[38;2;253;253;253mr[0m[38;2;242;242;242m2[0m[38;2;254;254;254mX[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255mr[0m[38;2;153;152;151mG[0m[38;2;29;29;30ms[0m[38;2;6;6;6m,[0m[38;2;52;52;56mA[0m[38;2;73;73;80m3[0m[38;2;78;79;86m3[0m[38;2;78;78;86m3[0m[38;2;77;77;84m3[0m[38;2;86;86;94mh[0m[38;2;86;87;95mh[0m[38;2;58;59;64m2[0m[38;2;1;1;1m.[0m[38;2;10;10;13m:[0m[38;2;13;14;20m;[0m[38;2;3;4;6m:[0m[38;2;0;0;0m.[0m[38;2;45;45;45m:[0m[38;2;108;108;108m:[0m[38;2;105;105;106m:[0m[38;2;104;104;104m:[0m[38;2;114;114;114m;[0m[38;2;135;135;135m:[0m[38;2;149;149;149mh[0m[38;2;119;119;120mS[0m[38;2;203;203;203m3[0m[38;2;222;222;222m,[0m[38;2;232;232;232m,[0m[38;2;244;244;244m.[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255mi[0m[38;2;243;243;243mh[0m[38;2;252;252;252mX[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m,[0m[38;2;253;253;253mi[0m[38;2;255;255;255m;[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m:[0m[38;2;248;248;248mH[0m[38;2;205;205;206mB[0m[38;2;195;195;196m&[0m[38;2;234;231;224m9[0m[38;2;255;232;184mB[0m[38;2;255;221;148m@[0m[38;2;242;209;142m&[0m[38;2;40;35;29mr[0m[38;2;140;131;77mG[0m[38;2;255;251;143m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;244;138m@[0m[38;2;255;246;139m@[0m[38;2;255;249;141m@[0m[38;2;255;252;143m@[0m[38;2;252;242;137m@[0m[38;2;201;193;110mB[0m[38;2;97;93;55m3[0m");
    $display("[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;254;254;253ms[0m[38;2;240;239;239mG[0m[38;2;211;210;212mB[0m[38;2;195;195;196m&[0m[38;2;213;212;213mB[0m[38;2;240;240;240mH[0m[38;2;255;255;255ms[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;254;254;254m3[0m[38;2;213;213;214m&[0m[38;2;191;191;193m&[0m[38;2;239;239;240m#[0m[38;2;255;255;255mr[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255ms[0m[38;2;235;234;235mB[0m[38;2;78;77;78m3[0m[38;2;15;15;16m:[0m[38;2;31;31;37mr[0m[38;2;39;39;48ms[0m[38;2;38;39;47ms[0m[38;2;37;38;46ms[0m[38;2;36;36;41ms[0m[38;2;31;31;35mr[0m[38;2;17;17;21m;[0m[38;2;13;13;18m:[0m[38;2;28;29;34mi[0m[38;2;38;38;42ms[0m[38;2;38;38;39ms[0m[38;2;11;11;12m,[0m[38;2;16;16;18m;[0m[38;2;17;17;20mi[0m[38;2;2;2;2m,[0m[38;2;8;8;8m:[0m[38;2;12;12;12m;[0m[38;2;4;3;4m:[0m[38;2;0;0;0m.[0m[38;2;3;2;2m.[0m[38;2;13;13;13m:[0m[38;2;26;25;26m;[0m[38;2;46;46;47mr[0m[38;2;84;84;85mA[0m[38;2;111;111;113mX[0m[38;2;135;135;135mi[0m[38;2;184;184;184m,[0m[38;2;235;235;235m.[0m[38;2;255;255;255mS[0m[38;2;180;180;181m&[0m[38;2;251;251;251mS[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;251;251;251m3[0m[38;2;219;219;219mB[0m[38;2;187;186;188m&[0m[38;2;219;219;220mB[0m[38;2;255;255;255m5[0m[38;2;255;253;244mi[0m[38;2;254;231;185m#[0m[38;2;255;220;146m@[0m[38;2;249;215;143m@[0m[38;2;54;47;36mX[0m[38;2;112;107;65mM[0m[38;2;255;250;142m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;252;143m@[0m[38;2;209;199;114mB[0m[38;2;77;72;43m2[0m");
    $display("[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m:[0m[38;2;249;249;249m5[0m[38;2;226;226;226m#[0m[38;2;200;200;202m&[0m[38;2;198;198;199m&[0m[38;2;216;215;216m#[0m[38;2;248;248;248mh[0m[38;2;255;255;255m;[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255ms[0m[38;2;235;235;235m#[0m[38;2;197;196;197m&[0m[38;2;203;203;204mB[0m[38;2;253;253;253mG[0m[38;2;255;255;255m:[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;249;249;249m [0m[38;2;156;155;155ms[0m[38;2;55;55;56mA[0m[38;2;16;17;22m;[0m[38;2;16;17;22m;[0m[38;2;24;24;31mi[0m[38;2;14;15;20m:[0m[38;2;4;4;7m.[0m[38;2;7;8;9m,[0m[38;2;34;34;36mr[0m[38;2;85;86;88mh[0m[38;2;152;154;157m9[0m[38;2;202;205;208m@[0m[38;2;219;222;226m@[0m[38;2;226;229;234m@[0m[38;2;195;197;202m&[0m[38;2;144;145;148m#[0m[38;2;119;120;123mG[0m[38;2;156;157;160m9[0m[38;2;205;207;211m@[0m[38;2;203;205;210m@[0m[38;2;179;181;184m&[0m[38;2;139;140;144m#[0m[38;2;91;91;93mh[0m[38;2;47;47;48mX[0m[38;2;20;20;22m;[0m[38;2;15;15;16m:[0m[38;2;31;30;32mr[0m[38;2;71;71;74m3[0m[38;2;114;114;117mS[0m[38;2;115;115;119mG[0m[38;2;95;95;96m5[0m[38;2;101;100;98m3[0m[38;2;145;144;144m#[0m[38;2;250;250;249m2[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;254m [0m[38;2;243;243;243mS[0m[38;2;212;212;212m9[0m[38;2;249;249;249mM[0m[38;2;255;255;255m,[0m[38;2;255;255;255m [0m[38;2;255;251;242mr[0m[38;2;254;232;187m#[0m[38;2;255;219;146m@[0m[38;2;253;219;145m@[0m[38;2;66;59;38mA[0m[38;2;101;96;58mh[0m[38;2;255;250;142m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;252;143m@[0m[38;2;198;189;108mB[0m[38;2;36;34;21mr[0m[38;2;130;118;89mh[0m");
    $display("[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255mr[0m[38;2;239;239;239mG[0m[38;2;198;198;199mB[0m[38;2;176;175;176m&[0m[38;2;193;192;193mB[0m[38;2;231;231;231mS[0m[38;2;252;252;251m2[0m[38;2;254;255;255m.[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m.[0m[38;2;181;180;180m3[0m[38;2;31;31;31ms[0m[38;2;74;73;74m3[0m[38;2;205;204;205m9[0m[38;2;255;255;255mh[0m[38;2;255;255;255m.[0m[38;2;255;255;255m [0m[38;2;231;231;231m:[0m[38;2;54;54;54m;[0m[38;2;2;2;3m.[0m[38;2;16;16;20m:[0m[38;2;13;14;19m:[0m[38;2;17;18;22m;[0m[38;2;51;52;55mA[0m[38;2;112;113;116mG[0m[38;2;175;177;182mB[0m[38;2;220;222;227m@[0m[38;2;241;244;249m@[0m[38;2;243;246;252m@[0m[38;2;239;242;248m@[0m[38;2;238;241;246m@[0m[38;2;237;240;245m@[0m[38;2;240;243;248m@[0m[38;2;243;246;251m@[0m[38;2;243;246;252m@[0m[38;2;243;246;251m@[0m[38;2;239;242;247m@[0m[38;2;239;242;247m@[0m[38;2;242;245;250m@[0m[38;2;244;247;252m@[0m[38;2;241;245;250m@[0m[38;2;223;226;231m@[0m[38;2;180;182;186m&[0m[38;2;121;122;125mS[0m[38;2;55;54;57mA[0m[38;2;15;15;16m:[0m[38;2;18;17;19m:[0m[38;2;66;66;68m2[0m[38;2;139;140;144m#[0m[38;2;163;165;169mB[0m[38;2;113;113;115mG[0m[38;2;87;87;87ms[0m[38;2;145;145;145m,[0m[38;2;228;228;228m.[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m.[0m[38;2;255;255;255m5[0m[38;2;246;246;246mh[0m[38;2;255;255;255mi[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255mi[0m[38;2;236;236;237mS[0m[38;2;224;225;225m#[0m[38;2;254;254;254m2[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;252;246mi[0m[38;2;254;233;190m#[0m[38;2;255;220;147m@[0m[38;2;255;221;146m@[0m[38;2;71;63;41mA[0m[38;2;97;93;55m3[0m[38;2;255;249;141m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;252;143m@[0m[38;2;197;188;108mB[0m[38;2;33;31;19mr[0m[38;2;144;129;94mM[0m[38;2;255;246;215mM[0m");
    $display("[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m:[0m[38;2;250;250;250m3[0m[38;2;219;219;219m9[0m[38;2;172;172;173mB[0m[38;2;223;223;223m&[0m[38;2;254;254;254mi[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;227;227;227m:[0m[38;2;33;33;33m:[0m[38;2;40;40;44ms[0m[38;2;42;42;46ms[0m[38;2;20;20;21mi[0m[38;2;134;134;134mS[0m[38;2;240;240;240m9[0m[38;2;255;255;255mA[0m[38;2;229;229;228m.[0m[38;2;89;89;89m;[0m[38;2;13;13;14m:[0m[38;2;36;36;37mr[0m[38;2;100;101;103mM[0m[38;2;170;172;176mB[0m[38;2;214;217;221m@[0m[38;2;245;248;253m@[0m[38;2;242;245;250m@[0m[38;2;238;241;246m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;239;242;247m@[0m[38;2;224;227;231m@[0m[38;2;186;188;192m&[0m[38;2;205;207;211m@[0m[38;2;176;177;181mB[0m[38;2;82;82;85m3[0m[38;2;26;27;29mi[0m[38;2;19;19;21m;[0m[38;2;63;63;65m2[0m[38;2;176;178;182m&[0m[38;2;212;215;220m@[0m[38;2;133;134;137m#[0m[38;2;79;79;80m2[0m[38;2;142;142;142m:[0m[38;2;237;237;237m.[0m[38;2;255;255;255m [0m[38;2;255;255;255m.[0m[38;2;224;224;224mh[0m[38;2;129;129;129mS[0m[38;2;69;68;69m5[0m[38;2;89;89;87mr[0m[38;2;183;183;184m:[0m[38;2;255;255;255m.[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;253;253;253m5[0m[38;2;212;212;213m9[0m[38;2;228;228;229m9[0m[38;2;255;255;255ms[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;253;249m;[0m[38;2;254;234;193mS[0m[38;2;255;220;148m@[0m[38;2;254;220;145m@[0m[38;2;69;61;40mA[0m[38;2;97;93;55m3[0m[38;2;255;249;141m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;252;143m@[0m[38;2;192;183;106m9[0m[38;2;34;31;20mr[0m[38;2;147;130;92mG[0m[38;2;255;244;208mG[0m[38;2;255;254;251m:[0m");
    $display("[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m.[0m[38;2;255;255;255m;[0m[38;2;253;253;253m;[0m[38;2;255;255;254m.[0m[38;2;253;253;253m3[0m[38;2;223;223;224m#[0m[38;2;235;235;235mG[0m[38;2;253;253;253mX[0m[38;2;255;255;255m.[0m[38;2;255;255;255m [0m[38;2;255;255;255m.[0m[38;2;109;109;109mi[0m[38;2;13;13;15m;[0m[38;2;81;81;89mh[0m[38;2;86;86;94mh[0m[38;2;61;62;67m2[0m[38;2;11;11;12m:[0m[38;2;76;76;77m3[0m[38;2;130;130;131mG[0m[38;2;47;47;48mi[0m[38;2;33;33;36ms[0m[38;2;100;100;103mM[0m[38;2;201;204;208m@[0m[38;2;192;194;198m&[0m[38;2;154;155;159m9[0m[38;2;217;220;225m@[0m[38;2;237;240;245m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;236;239;244m@[0m[38;2;191;193;197m&[0m[38;2;91;91;93mh[0m[38;2;137;138;142m#[0m[38;2;237;240;246m@[0m[38;2;191;193;197m&[0m[38;2;108;109;112mH[0m[38;2;47;47;50mX[0m[38;2;17;17;19m:[0m[38;2;114;115;118mG[0m[38;2;240;244;249m@[0m[38;2;230;233;238m@[0m[38;2;169;171;175m&[0m[38;2;104;104;106m5[0m[38;2;142;142;142m:[0m[38;2;106;106;107m;[0m[38;2;49;49;51mX[0m[38;2;44;44;49mX[0m[38;2;66;66;73m5[0m[38;2;37;37;41mX[0m[38;2;29;29;29m;[0m[38;2;230;230;230m:[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;254;254;254m,[0m[38;2;252;252;252mX[0m[38;2;246;246;247m2[0m[38;2;255;255;255m;[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;253;250m:[0m[38;2;254;235;196mG[0m[38;2;255;220;150m@[0m[38;2;254;219;144m@[0m[38;2;65;58;38mA[0m[38;2;101;96;57mh[0m[38;2;255;250;142m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;252;143m@[0m[38;2;186;177;102m9[0m[38;2;33;29;20mi[0m[38;2;154;134;94mG[0m[38;2;255;242;199mS[0m[38;2;255;253;247m;[0m[38;2;255;255;255m [0m");
    $display("[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;254;254;254mX[0m[38;2;234;234;234m#[0m[38;2;204;203;204m&[0m[38;2;198;198;200m&[0m[38;2;219;219;220m9[0m[38;2;250;250;250mh[0m[38;2;202;202;201mr[0m[38;2;16;16;16m:[0m[38;2;59;60;65m2[0m[38;2;85;85;93mh[0m[38;2;83;83;91mh[0m[38;2;86;86;94mh[0m[38;2;72;72;79m5[0m[38;2;10;11;12m,[0m[38;2;0;0;0m.[0m[38;2;49;49;53mA[0m[38;2;159;161;165mB[0m[38;2;235;237;241m@[0m[38;2;118;119;122mG[0m[38;2;91;91;94mM[0m[38;2;219;222;227m@[0m[38;2;239;242;247m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;236;239;244m@[0m[38;2;236;239;244m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;241;244;249m@[0m[38;2;227;229;234m@[0m[38;2;86;87;88mh[0m[38;2;93;94;97mM[0m[38;2;241;244;250m@[0m[38;2;242;245;250m@[0m[38;2;187;188;193m&[0m[38;2;63;63;66m2[0m[38;2;6;6;8m,[0m[38;2;103;103;106mH[0m[38;2;213;216;220m@[0m[38;2;140;141;144m#[0m[38;2;57;57;58m2[0m[38;2;38;38;42mX[0m[38;2;64;64;71m5[0m[38;2;80;80;88mh[0m[38;2;85;85;93mh[0m[38;2;85;85;94mh[0m[38;2;71;71;77m5[0m[38;2;7;7;8m:[0m[38;2;179;179;179m;[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;254;253;253mA[0m[38;2;213;213;214m&[0m[38;2;222;222;222m&[0m[38;2;254;254;254mX[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;254;250m:[0m[38;2;253;235;198m9[0m[38;2;254;219;147m@[0m[38;2;253;220;145m@[0m[38;2;59;53;36mX[0m[38;2;73;69;40m2[0m[38;2;255;247;140m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;245;139m@[0m[38;2;255;253;144m@[0m[38;2;174;166;96m#[0m[38;2;31;29;19mi[0m[38;2;164;143;97mS[0m[38;2;255;240;190m#[0m[38;2;255;254;244mr[0m[38;2;255;255;255m,[0m[38;2;254;254;254m,[0m");
    $display("[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;254;254;254m;[0m[38;2;243;243;244m5[0m[38;2;249;249;249mA[0m[38;2;255;255;255m;[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255mi[0m[38;2;246;246;246mh[0m[38;2;219;219;219m9[0m[38;2;198;198;199m&[0m[38;2;65;64;63mA[0m[38;2;23;23;25mi[0m[38;2;80;80;88m3[0m[38;2;79;79;87m3[0m[38;2;76;77;85m3[0m[38;2;74;75;82m3[0m[38;2;77;77;85m3[0m[38;2;41;42;46ms[0m[38;2;40;40;41ms[0m[38;2;186;188;192m&[0m[38;2;229;230;236m@[0m[38;2;87;87;89mh[0m[38;2;83;84;86mh[0m[38;2;226;228;233m@[0m[38;2;239;242;247m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;238;241;246m@[0m[38;2;237;240;245m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;236;239;244m@[0m[38;2;228;231;235m@[0m[38;2;233;236;241m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;240;243;248m@[0m[38;2;218;220;225m@[0m[38;2;35;35;36mr[0m[38;2;136;137;141m#[0m[38;2;243;246;252m@[0m[38;2;245;248;253m@[0m[38;2;176;177;180mB[0m[38;2;23;22;23m;[0m[38;2;5;5;5m.[0m[38;2;27;27;28mi[0m[38;2;39;38;43ms[0m[38;2;70;70;77m5[0m[38;2;85;85;93mh[0m[38;2;83;83;91mh[0m[38;2;83;82;90mh[0m[38;2;83;83;90mh[0m[38;2;84;84;92mh[0m[38;2;76;77;84m3[0m[38;2;9;9;10m;[0m[38;2;155;155;155m;[0m[38;2;255;255;255mi[0m[38;2;239;239;239mG[0m[38;2;224;224;225m#[0m[38;2;253;252;252m5[0m[38;2;252;252;252mi[0m[38;2;255;255;255m;[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m,[0m[38;2;252;252;252mA[0m[38;2;233;233;233mG[0m[38;2;217;216;217m9[0m[38;2;252;251;249mG[0m[38;2;254;236;200mS[0m[38;2;254;220;150m@[0m[38;2;254;219;145m@[0m[38;2;59;54;36mX[0m[38;2;54;52;32mX[0m[38;2;254;243;138m@[0m[38;2;255;244;139m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;246;140m@[0m[38;2;251;242;138m@[0m[38;2;142;135;78mG[0m[38;2;30;27;19mi[0m[38;2;173;151;99m#[0m[38;2;255;234;178m&[0m[38;2;243;236;221mS[0m[38;2;227;227;228m#[0m[38;2;211;211;212mB[0m[38;2;211;211;211mB[0m");
    $display("[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;254;254;253mX[0m[38;2;225;225;225mB[0m[38;2;201;201;202m&[0m[38;2;205;205;206m&[0m[38;2;218;218;218m9[0m[38;2;235;234;234mH[0m[38;2;249;249;249m2[0m[38;2;254;254;254m,[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m.[0m[38;2;175;175;175mA[0m[38;2;3;3;3m,[0m[38;2;30;31;38mr[0m[38;2;38;39;49ms[0m[38;2;37;38;48ms[0m[38;2;35;36;47ms[0m[38;2;34;35;45ms[0m[38;2;18;19;24m;[0m[38;2;58;58;60mA[0m[38;2;218;221;224m@[0m[38;2;227;230;238m@[0m[38;2;80;81;87m3[0m[38;2;91;91;93mh[0m[38;2;231;234;239m@[0m[38;2;239;242;247m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;240;243;248m@[0m[38;2;210;213;218m@[0m[38;2;204;206;211m@[0m[38;2;238;241;246m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;242;245;250m@[0m[38;2;149;150;154m9[0m[38;2;165;167;171mB[0m[38;2;241;244;249m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;233;236;241m@[0m[38;2;237;240;245m@[0m[38;2;245;249;254m@[0m[38;2;140;142;145m#[0m[38;2;35;35;36mr[0m[38;2;221;224;228m@[0m[38;2;239;242;247m@[0m[38;2;243;246;251m@[0m[38;2;100;101;103mH[0m[38;2;0;0;0m [0m[38;2;6;6;7m,[0m[38;2;37;38;45ms[0m[38;2;42;43;53mX[0m[38;2;41;42;52mX[0m[38;2;43;44;52mX[0m[38;2;44;45;53mX[0m[38;2;45;45;54mX[0m[38;2;46;47;56mX[0m[38;2;44;44;52mX[0m[38;2;5;5;6m,[0m[38;2;154;153;151mh[0m[38;2;217;217;217m&[0m[38;2;188;187;188m&[0m[38;2;231;231;232mB[0m[38;2;255;255;254mr[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m.[0m[38;2;254;253;253ms[0m[38;2;240;241;241mH[0m[38;2;216;215;216mB[0m[38;2;197;197;198m&[0m[38;2;207;207;207mB[0m[38;2;233;234;234mS[0m[38;2;254;254;253mA[0m[38;2;255;237;203mH[0m[38;2;254;220;151m&[0m[38;2;255;225;149m@[0m[38;2;97;86;57m3[0m[38;2;68;64;39mA[0m[38;2;255;246;139m@[0m[38;2;255;244;138m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;247;140m@[0m[38;2;245;236;135m@[0m[38;2;86;81;48m5[0m[38;2;23;20;14m;[0m[38;2;189;164;111m9[0m[38;2;255;234;177m&[0m[38;2;227;218;203mB[0m[38;2;210;210;211mB[0m[38;2;220;220;221m#[0m[38;2;236;236;236mM[0m[38;2;249;249;249m2[0m");
    $display("[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m,[0m[38;2;254;254;253mr[0m[38;2;244;244;244m3[0m[38;2;229;228;229mS[0m[38;2;211;211;212m9[0m[38;2;230;230;230m9[0m[38;2;255;255;255mr[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;254;254;254m.[0m[38;2;255;255;255m,[0m[38;2;255;255;255m.[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;254;254;254m.[0m[38;2;80;80;80m;[0m[38;2;0;0;0m,[0m[38;2;19;20;27mi[0m[38;2;20;21;27m;[0m[38;2;19;20;25m;[0m[38;2;19;20;24m;[0m[38;2;13;13;16m:[0m[38;2;8;7;7m,[0m[38;2;183;185;188m&[0m[38;2;233;238;246m@[0m[38;2;89;94;104mM[0m[38;2;31;31;32mr[0m[38;2;224;226;231m@[0m[38;2;239;242;248m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;238;241;247m@[0m[38;2;211;214;217m@[0m[38;2;58;57;59mA[0m[38;2;183;185;190m&[0m[38;2;241;244;249m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;243;247;252m@[0m[38;2;104;104;106mH[0m[38;2;77;77;79m3[0m[38;2;243;246;251m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;236;239;244m@[0m[38;2;212;214;218m@[0m[38;2;238;241;246m@[0m[38;2;210;212;217m@[0m[38;2;25;25;26mi[0m[38;2;165;165;169mB[0m[38;2;242;245;250m@[0m[38;2;233;235;237m@[0m[38;2;190;191;193m&[0m[38;2;23;21;20m;[0m[38;2;24;23;23m;[0m[38;2;8;8;10m,[0m[38;2;22;23;30mi[0m[38;2;23;24;31mi[0m[38;2;26;26;35mi[0m[38;2;28;29;38mr[0m[38;2;26;27;37mi[0m[38;2;28;29;39mr[0m[38;2;20;21;27m;[0m[38;2;0;0;0m.[0m[38;2;140;140;141m9[0m[38;2;223;223;224mB[0m[38;2;253;253;253m3[0m[38;2;255;255;255m.[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;254;254;254mX[0m[38;2;220;220;220m&[0m[38;2;197;196;197m&[0m[38;2;224;223;224m#[0m[38;2;249;249;249m3[0m[38;2;255;255;255m;[0m[38;2;255;255;255m [0m[38;2;255;251;242mi[0m[38;2;255;233;187m#[0m[38;2;255;226;155m@[0m[38;2;255;232;154m@[0m[38;2;93;80;55m3[0m[38;2;93;88;52m3[0m[38;2;255;251;143m@[0m[38;2;255;250;142m@[0m[38;2;255;249;141m@[0m[38;2;255;247;138m@[0m[38;2;255;250;141m@[0m[38;2;255;251;142m@[0m[38;2;255;251;142m@[0m[38;2;255;250;142m@[0m[38;2;249;241;137m@[0m[38;2;91;87;52m3[0m[38;2;62;54;38mA[0m[38;2;220;193;130mB[0m[38;2;255;236;185m9[0m[38;2;255;248;234mA[0m[38;2;255;255;255m:[0m[38;2;255;255;255m,[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m");
    $display("[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m.[0m[38;2;255;255;255m.[0m[38;2;255;255;255m.[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;252;252;252mh[0m[38;2;215;215;215mB[0m[38;2;214;214;214m9[0m[38;2;242;242;242mG[0m[38;2;254;254;254m:[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;210;210;210m,[0m[38;2;166;166;166m:[0m[38;2;73;73;73m;[0m[38;2;0;0;0m.[0m[38;2;14;14;17m:[0m[38;2;14;16;21m:[0m[38;2;10;13;22m:[0m[38;2;17;18;22m;[0m[38;2;120;123;129mS[0m[38;2;125;135;154m#[0m[38;2;3;4;7m.[0m[38;2;112;113;115mG[0m[38;2;244;247;252m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;242;245;250m@[0m[38;2;114;115;117mG[0m[38;2;46;46;48mX[0m[38;2;228;231;236m@[0m[38;2;237;240;245m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;243;246;252m@[0m[38;2;117;118;120mG[0m[38;2;18;18;19m;[0m[38;2;191;193;197m&[0m[38;2;240;243;248m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;242;245;250m@[0m[38;2;131;132;134mS[0m[38;2;165;167;170mB[0m[38;2;239;242;247m@[0m[38;2;57;57;59mA[0m[38;2;51;51;52mX[0m[38;2;73;74;79m3[0m[38;2;57;65;88m5[0m[38;2;55;63;88m5[0m[38;2;24;30;49mr[0m[38;2;10;11;13m,[0m[38;2;1;1;0m [0m[38;2;13;14;17m:[0m[38;2;17;17;21m;[0m[38;2;13;13;16m:[0m[38;2;7;8;9m,[0m[38;2;41;41;45ms[0m[38;2;16;16;19m:[0m[38;2;20;20;22m;[0m[38;2;122;122;123mM[0m[38;2;245;244;245mH[0m[38;2;255;255;255m;[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m.[0m[38;2;255;255;255ms[0m[38;2;232;232;232mS[0m[38;2;235;235;236mS[0m[38;2;255;255;255mi[0m[38;2;254;254;254m,[0m[38;2;251;251;251mr[0m[38;2;255;255;255mi[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;254m.[0m[38;2;255;251;230m5[0m[38;2;255;232;181m9[0m[38;2;190;165;114m9[0m[38;2;131;115;80mH[0m[38;2;48;42;31ms[0m[38;2;177;168;96m9[0m[38;2;246;238;136m@[0m[38;2;108;102;58mh[0m[38;2;114;108;68mM[0m[38;2;167;158;111m#[0m[38;2;153;146;91mS[0m[38;2;161;152;88m#[0m[38;2;170;162;90m#[0m[38;2;204;198;112mB[0m[38;2;119;112;66mM[0m[38;2;55;48;35mX[0m[38;2;233;203;135m&[0m[38;2;255;231;171m&[0m[38;2;255;246;227m2[0m[38;2;255;255;255m.[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m");
    $display("[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;254;254;254m;[0m[38;2;246;246;246m5[0m[38;2;232;232;232mM[0m[38;2;241;241;241mH[0m[38;2;254;254;254m:[0m[38;2;255;255;255m [0m[38;2;253;252;252m2[0m[38;2;239;237;237mM[0m[38;2;247;246;245m5[0m[38;2;255;255;255mi[0m[38;2;255;255;255m,[0m[38;2;161;161;160m;[0m[38;2;23;22;19m,[0m[38;2;17;24;45mi[0m[38;2;52;80;159mM[0m[38;2;51;77;153mM[0m[38;2;10;14;25m:[0m[38;2;72;80;91m3[0m[38;2;48;53;63mA[0m[38;2;2;2;1m.[0m[38;2;176;178;182m&[0m[38;2;242;245;250m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;236;239;244m@[0m[38;2;233;235;240m@[0m[38;2;49;48;50mX[0m[38;2;117;117;120mG[0m[38;2;243;246;252m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;243;246;251m@[0m[38;2;127;127;130mS[0m[38;2;0;0;0m [0m[38;2;67;67;69m5[0m[38;2;234;237;242m@[0m[38;2;236;239;244m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;243;246;252m@[0m[38;2;125;126;128mS[0m[38;2;75;75;76m3[0m[38;2;234;236;241m@[0m[38;2;71;70;68m5[0m[38;2;19;17;14m:[0m[38;2;7;7;9m,[0m[38;2;44;69;144mh[0m[38;2;53;84;175mH[0m[38;2;47;71;142mh[0m[38;2;6;6;8m,[0m[38;2;3;1;0m.[0m[38;2;13;13;15m:[0m[38;2;33;34;45mr[0m[38;2;24;25;32mi[0m[38;2;9;9;9m,[0m[38;2;185;186;190m&[0m[38;2;120;121;124mS[0m[38;2;49;49;49mr[0m[38;2;252;252;252ms[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m.[0m[38;2;255;254;254mX[0m[38;2;237;237;237mG[0m[38;2;212;211;211m9[0m[38;2;239;239;239m&[0m[38;2;226;226;226m#[0m[38;2;237;237;237mG[0m[38;2;254;254;254m;[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m.[0m[38;2;206;202;190mA[0m[38;2;83;78;66mA[0m[38;2;83;78;75m3[0m[38;2;175;163;161mB[0m[38;2;95;89;73mh[0m[38;2;239;227;128m&[0m[38;2;130;122;70mH[0m[38;2;31;29;34mr[0m[38;2;162;149;146m9[0m[38;2;201;189;184m&[0m[38;2;172;160;157mB[0m[38;2;136;128;127mS[0m[38;2;91;86;87mh[0m[38;2;41;38;35ms[0m[38;2;0;0;0m [0m[38;2;79;69;46m2[0m[38;2;242;210;144m&[0m[38;2;255;232;182m9[0m[38;2;255;249;237ms[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m");
    $display("[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;253;252;252mh[0m[38;2;222;222;223mB[0m[38;2;204;204;205m&[0m[38;2;206;206;207m&[0m[38;2;185;185;185m#[0m[38;2;102;104;113mr[0m[38;2;56;64;88mX[0m[38;2;31;46;89mA[0m[38;2;56;88;178mH[0m[38;2;43;67;135m3[0m[38;2;16;22;41mi[0m[38;2;32;40;59ms[0m[38;2;2;2;2m.[0m[38;2;17;17;18m:[0m[38;2;206;208;214m@[0m[38;2;239;242;247m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;240;243;248m@[0m[38;2;195;197;202m&[0m[38;2;14;14;14m:[0m[38;2;155;156;159m9[0m[38;2;245;248;254m@[0m[38;2;236;239;244m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;243;246;251m@[0m[38;2;130;130;133mS[0m[38;2;10;9;6m,[0m[38;2;19;19;17m;[0m[38;2;190;192;196m&[0m[38;2;240;244;249m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;242;245;251m@[0m[38;2;154;155;158m9[0m[38;2;31;30;31mr[0m[38;2;54;54;57mA[0m[38;2;30;38;64ms[0m[38;2;27;39;74mX[0m[38;2;29;43;83mA[0m[38;2;52;80;161mM[0m[38;2;57;88;179mH[0m[38;2;36;54;106m2[0m[38;2;14;19;35m;[0m[38;2;19;26;48mr[0m[38;2;8;11;17m,[0m[38;2;10;10;11m,[0m[38;2;16;16;21m:[0m[38;2;25;24;25m;[0m[38;2;219;221;226m@[0m[38;2;192;194;198m&[0m[38;2;33;32;32m;[0m[38;2;225;225;225m,[0m[38;2;255;255;255mr[0m[38;2;243;243;243mM[0m[38;2;220;220;220m9[0m[38;2;198;198;200m&[0m[38;2;204;204;205m&[0m[38;2;229;229;229m#[0m[38;2;250;250;250m5[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m,[0m[38;2;242;241;239m;[0m[38;2;238;238;239m2[0m[38;2;153;153;152mX[0m[38;2;41;40;41mr[0m[38;2;154;144;139m9[0m[38;2;252;237;226m@[0m[38;2;247;229;221m@[0m[38;2;91;86;68m3[0m[38;2;148;140;76mG[0m[38;2;13;13;8m,[0m[38;2;77;74;73m5[0m[38;2;138;129;124mS[0m[38;2;180;168;160mB[0m[38;2;228;212;203m@[0m[38;2;251;234;223m@[0m[38;2;255;241;230m@[0m[38;2;231;215;206m@[0m[38;2;169;160;153m9[0m[38;2;54;51;51mA[0m[38;2;71;62;44mA[0m[38;2;248;228;181m#[0m[38;2;255;251;239ms[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m");
    $display("[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m.[0m[38;2;255;255;255mi[0m[38;2;250;250;250m5[0m[38;2;167;166;163m3[0m[38;2;4;12;34mr[0m[38;2;38;61;128m3[0m[38;2;43;65;127m3[0m[38;2;55;84;171mH[0m[38;2;53;82;166mM[0m[38;2;34;50;97m2[0m[38;2;28;39;71mX[0m[38;2;0;0;0m [0m[38;2;28;28;30mi[0m[38;2;221;223;228m@[0m[38;2;239;242;247m@[0m[38;2;237;240;244m@[0m[38;2;237;240;245m@[0m[38;2;240;243;248m@[0m[38;2;91;91;93mh[0m[38;2;0;0;0m [0m[38;2;167;168;171mB[0m[38;2;228;231;235m@[0m[38;2;232;235;240m@[0m[38;2;237;240;245m@[0m[38;2;237;240;245m@[0m[38;2;237;240;245m@[0m[38;2;237;240;245m@[0m[38;2;237;240;246m@[0m[38;2;238;241;246m@[0m[38;2;245;248;253m@[0m[38;2;141;142;146m#[0m[38;2;46;36;28mr[0m[38;2;43;33;27mr[0m[38;2;118;120;123mG[0m[38;2;249;252;255m@[0m[38;2;243;246;251m@[0m[38;2;243;246;251m@[0m[38;2;244;247;252m@[0m[38;2;250;254;255m@[0m[38;2;185;186;191m&[0m[38;2;56;55;55mA[0m[38;2;4;5;9m.[0m[38;2;42;64;129m3[0m[38;2;44;68;135m3[0m[38;2;43;65;131m3[0m[38;2;53;81;162mM[0m[38;2;55;86;173mH[0m[38;2;54;84;169mH[0m[38;2;56;87;175mH[0m[38;2;55;85;170mH[0m[38;2;15;20;36m;[0m[38;2;0;0;0m [0m[38;2;0;0;3m.[0m[38;2;43;43;44ms[0m[38;2;230;233;237m@[0m[38;2;222;224;230m@[0m[38;2;52;52;53mX[0m[38;2;185;183;182m#[0m[38;2;186;185;186m&[0m[38;2;191;191;191m&[0m[38;2;222;222;222m9[0m[38;2;246;246;246mh[0m[38;2;255;255;255mi[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m.[0m[38;2;255;255;255m;[0m[38;2;255;255;255mX[0m[38;2;233;233;233m3[0m[38;2;182;183;183m3[0m[38;2;105;104;105mA[0m[38;2;37;35;34m;[0m[38;2;28;28;29mr[0m[38;2;11;11;11m;[0m[38;2;180;167;160mB[0m[38;2;255;246;235m@[0m[38;2;255;243;231m@[0m[38;2;213;198;190m&[0m[38;2;28;26;26mi[0m[38;2;92;86;83mh[0m[38;2;186;175;168mB[0m[38;2;234;218;208m@[0m[38;2;252;234;223m@[0m[38;2;254;236;225m@[0m[38;2;249;231;220m@[0m[38;2;248;230;220m@[0m[38;2;252;234;223m@[0m[38;2;255;242;231m@[0m[38;2;255;253;241m@[0m[38;2;102;95;92mM[0m[38;2;61;58;52ms[0m[38;2;249;240;216mh[0m[38;2;255;255;252m:[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m");
    $display("[38;2;223;222;223mG[0m[38;2;231;231;231mH[0m[38;2;237;237;237m3[0m[38;2;245;245;244m2[0m[38;2;249;249;249ms[0m[38;2;254;254;254mi[0m[38;2;255;255;255m:[0m[38;2;255;255;255m.[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;246;246;246m [0m[38;2;171;171;171m:[0m[38;2;73;72;69m:[0m[38;2;7;12;28m;[0m[38;2;47;76;158mM[0m[38;2;45;70;143mh[0m[38;2;5;6;9m,[0m[38;2;2;2;0m.[0m[38;2;16;13;11m:[0m[38;2;73;69;68m5[0m[38;2;229;232;237m@[0m[38;2;229;232;238m@[0m[38;2;226;229;235m@[0m[38;2;227;231;236m@[0m[38;2;226;229;234m@[0m[38;2;59;59;61m2[0m[38;2;3;2;2m.[0m[38;2;94;94;97mM[0m[38;2;32;32;34mr[0m[38;2;103;105;107mH[0m[38;2;228;231;236m@[0m[38;2;222;225;230m@[0m[38;2;219;223;228m@[0m[38;2;217;220;225m@[0m[38;2;213;216;221m@[0m[38;2;211;214;219m@[0m[38;2;220;223;229m@[0m[38;2;178;181;185m&[0m[38;2;135;104;97mG[0m[38;2;151;122;114mS[0m[38;2;57;60;62m2[0m[38;2;179;180;185m&[0m[38;2;164;166;170mB[0m[38;2;154;156;160m9[0m[38;2;148;150;153m9[0m[38;2;124;125;129mS[0m[38;2;67;67;69m5[0m[38;2;49;47;47ms[0m[38;2;17;16;16m:[0m[38;2;5;5;5m.[0m[38;2;23;21;20m;[0m[38;2;12;14;24m:[0m[38;2;50;76;155mM[0m[38;2;56;88;182mH[0m[38;2;47;69;132m3[0m[38;2;23;31;55mr[0m[38;2;23;33;65ms[0m[38;2;1;1;1m.[0m[38;2;76;76;79m3[0m[38;2;89;90;92mh[0m[38;2;154;155;159m9[0m[38;2;242;245;250m@[0m[38;2;206;208;212m@[0m[38;2;34;34;35mr[0m[38;2;175;175;175mS[0m[38;2;241;242;242mG[0m[38;2;252;252;251mA[0m[38;2;255;255;255m.[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m.[0m[38;2;252;252;252m.[0m[38;2;218;218;218m.[0m[38;2;178;178;178m;[0m[38;2;138;137;138mM[0m[38;2;97;97;98mh[0m[38;2;87;87;88mM[0m[38;2;109;109;111mG[0m[38;2;141;141;142m9[0m[38;2;63;63;65m2[0m[38;2;31;28;27mi[0m[38;2;176;165;157mB[0m[38;2;255;247;236m@[0m[38;2;255;242;231m@[0m[38;2;226;211;202m@[0m[38;2;44;42;42ms[0m[38;2;62;58;56mA[0m[38;2;153;143;137m#[0m[38;2;139;130;125mS[0m[38;2;132;124;120mS[0m[38;2;150;140;134m#[0m[38;2;188;175;168mB[0m[38;2;217;203;194m@[0m[38;2;236;220;210m@[0m[38;2;224;207;198m@[0m[38;2;154;145;140m9[0m[38;2;203;189;182m&[0m[38;2;28;26;26mr[0m[38;2;156;147;128m5[0m[38;2;255;255;248mX[0m[38;2;255;255;255m.[0m[38;2;254;254;254m.[0m[38;2;255;255;255m [0m[38;2;255;255;255m.[0m[38;2;249;249;249m2[0m[38;2;233;232;232m3[0m[38;2;231;231;232mH[0m");
    $display("[38;2;225;225;225mG[0m[38;2;217;218;218m#[0m[38;2;212;211;211m9[0m[38;2;206;206;207mB[0m[38;2;206;206;206mB[0m[38;2;204;203;204mB[0m[38;2;210;210;210mB[0m[38;2;211;211;211m9[0m[38;2;219;219;219m#[0m[38;2;226;226;226mG[0m[38;2;232;231;231mM[0m[38;2;239;239;239m3[0m[38;2;246;246;246mA[0m[38;2;254;254;254m:[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;235;235;234m,[0m[38;2;138;138;137m:[0m[38;2;18;18;17m,[0m[38;2;39;42;52mX[0m[38;2;59;67;87m5[0m[38;2;47;54;73mA[0m[38;2;31;34;40mr[0m[38;2;12;14;18m:[0m[38;2;43;34;30mr[0m[38;2;108;96;91mM[0m[38;2;69;72;76m5[0m[38;2;60;61;65m2[0m[38;2;82;82;84m3[0m[38;2;121;117;116mG[0m[38;2;193;184;179m&[0m[38;2;201;185;179m&[0m[38;2;183;164;156mB[0m[38;2;115;109;104mH[0m[38;2;114;106;102mH[0m[38;2;126;118;113mG[0m[38;2;115;111;109mG[0m[38;2;106;103;102mH[0m[38;2;107;102;101mH[0m[38;2;107;102;100mH[0m[38;2;110;104;102mH[0m[38;2;114;109;107mH[0m[38;2;158;150;147m9[0m[38;2;215;204;197m@[0m[38;2;220;195;186m&[0m[38;2;197;182;175m&[0m[38;2;48;46;46mX[0m[38;2;0;0;0m [0m[38;2;0;0;0m [0m[38;2;0;0;0m [0m[38;2;0;0;0m [0m[38;2;15;13;12m:[0m[38;2;53;49;48mX[0m[38;2;155;146;139m9[0m[38;2;130;120;115mG[0m[38;2;4;5;6m.[0m[38;2;24;26;30mi[0m[38;2;23;28;45mr[0m[38;2;33;45;78mA[0m[38;2;35;46;77mA[0m[38;2;33;40;58ms[0m[38;2;12;11;7m,[0m[38;2;24;23;23m;[0m[38;2;59;60;62m2[0m[38;2;202;204;209m@[0m[38;2;229;232;237m@[0m[38;2;242;245;250m@[0m[38;2;242;246;251m@[0m[38;2;175;177;181m&[0m[38;2;33;33;33m;[0m[38;2;223;223;223m:[0m[38;2;151;151;151m,[0m[38;2;87;87;88mr[0m[38;2;87;87;87mi[0m[38;2;101;101;101m;[0m[38;2;117;117;117mr[0m[38;2;106;106;106m;[0m[38;2;73;73;74mi[0m[38;2;100;100;101mh[0m[38;2;146;146;147m9[0m[38;2;181;180;181m&[0m[38;2;211;211;212m@[0m[38;2;245;245;246m@[0m[38;2;255;255;255m@[0m[38;2;201;201;202m&[0m[38;2;30;29;30mi[0m[38;2;194;179;172m&[0m[38;2;255;247;235m@[0m[38;2;197;182;174m&[0m[38;2;86;81;78m3[0m[38;2;57;54;53mA[0m[38;2;72;68;65m5[0m[38;2;136;128;123mS[0m[38;2;172;161;154mB[0m[38;2;205;191;183m&[0m[38;2;233;217;207m@[0m[38;2;249;231;220m@[0m[38;2;255;237;226m@[0m[38;2;255;237;226m@[0m[38;2;255;237;226m@[0m[38;2;252;234;223m@[0m[38;2;229;217;208m@[0m[38;2;158;149;143m9[0m[38;2;15;15;15m:[0m[38;2;207;195;175m#[0m[38;2;217;215;210mB[0m[38;2;215;215;215mB[0m[38;2;252;252;253mM[0m[38;2;255;255;255m [0m[38;2;255;255;255m.[0m[38;2;243;243;243mS[0m[38;2;206;206;207m#[0m[38;2;224;224;224mS[0m");
    $display("[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m.[0m[38;2;255;255;255m,[0m[38;2;255;255;255m;[0m[38;2;251;251;251mr[0m[38;2;247;247;247mA[0m[38;2;240;240;240m5[0m[38;2;233;233;233mh[0m[38;2;228;228;228mH[0m[38;2;219;218;219mS[0m[38;2;216;216;217m#[0m[38;2;227;227;228m9[0m[38;2;254;254;254mX[0m[38;2;255;255;255m [0m[38;2;255;255;255m,[0m[38;2;244;244;244mG[0m[38;2;217;217;218mS[0m[38;2;233;233;233mG[0m[38;2;239;238;239mM[0m[38;2;219;218;218mX[0m[38;2;133;133;133m:[0m[38;2;74;74;75mX[0m[38;2;64;64;66m5[0m[38;2;15;15;16m:[0m[38;2;190;192;197m&[0m[38;2;230;233;239m@[0m[38;2;214;219;227m@[0m[38;2;202;208;219m@[0m[38;2;151;155;164m9[0m[38;2;13;13;14m:[0m[38;2;13;13;13m,[0m[38;2;39;37;36mi[0m[38;2;18;17;17m:[0m[38;2;17;16;16m:[0m[38;2;38;35;34mr[0m[38;2;72;67;64m5[0m[38;2;113;106;101mH[0m[38;2;155;145;139m9[0m[38;2;191;178;170m&[0m[38;2;226;211;201m@[0m[38;2;250;233;222m@[0m[38;2;251;232;221m@[0m[38;2;249;231;220m@[0m[38;2;250;232;221m@[0m[38;2;252;234;223m@[0m[38;2;255;237;226m@[0m[38;2;251;234;223m@[0m[38;2;166;155;149m9[0m[38;2;98;91;87mM[0m[38;2;44;42;40ms[0m[38;2;27;26;26mi[0m[38;2;43;41;40ms[0m[38;2;72;68;66m5[0m[38;2;115;108;104mH[0m[38;2;158;148;142m9[0m[38;2;190;176;169m&[0m[38;2;232;215;206m@[0m[38;2;253;236;225m@[0m[38;2;255;244;233m@[0m[38;2;76;71;68m5[0m[38;2;60;63;71m2[0m[38;2;168;177;194m&[0m[38;2;180;185;193m&[0m[38;2;195;196;198m&[0m[38;2;203;204;206m@[0m[38;2;199;200;202m&[0m[38;2;42;43;45ms[0m[38;2;19;20;22m;[0m[38;2;49;47;48mX[0m[38;2;26;26;27mi[0m[38;2;159;160;164mB[0m[38;2;244;247;252m@[0m[38;2;238;240;245m@[0m[38;2;81;81;83m3[0m[38;2;27;26;26m:[0m[38;2;62;62;63mi[0m[38;2;107;107;109mG[0m[38;2;225;225;226m@[0m[38;2;196;196;200m@[0m[38;2;116;114;122mS[0m[38;2;18;18;19mi[0m[38;2;69;69;72m3[0m[38;2;202;201;202m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;242;241;242m@[0m[38;2;50;50;52mX[0m[38;2;114;106;102mH[0m[38;2;255;242;230m@[0m[38;2;255;239;228m@[0m[38;2;108;102;99mH[0m[38;2;0;0;0m [0m[38;2;130;121;118mS[0m[38;2;255;242;231m@[0m[38;2;255;253;241m@[0m[38;2;255;250;238m@[0m[38;2;255;245;233m@[0m[38;2;255;240;229m@[0m[38;2;255;237;226m@[0m[38;2;254;236;225m@[0m[38;2;253;235;224m@[0m[38;2;253;235;224m@[0m[38;2;254;236;225m@[0m[38;2;255;243;231m@[0m[38;2;102;96;93mM[0m[38;2;67;63;55ms[0m[38;2;252;242;220mG[0m[38;2;245;244;242m5[0m[38;2;248;247;247m2[0m[38;2;254;254;254mi[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m");
    $display("[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m.[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m.[0m[38;2;255;255;255m2[0m[38;2;221;221;221mM[0m[38;2;155;155;155mG[0m[38;2;73;73;74m3[0m[38;2;72;71;72m3[0m[38;2;133;134;137m#[0m[38;2;215;218;224m@[0m[38;2;89;90;94mh[0m[38;2;58;58;60mA[0m[38;2;236;239;244m@[0m[38;2;238;241;246m@[0m[38;2;238;241;245m@[0m[38;2;240;242;247m@[0m[38;2;246;249;253m@[0m[38;2;119;121;126mS[0m[38;2;6;6;6m.[0m[38;2;159;150;144m#[0m[38;2;225;213;204m@[0m[38;2;188;175;167mB[0m[38;2;151;141;135m#[0m[38;2;116;108;103mH[0m[38;2;87;81;77m3[0m[38;2;69;64;62m2[0m[38;2;48;44;43mX[0m[38;2;14;14;13m:[0m[38;2;30;28;27mi[0m[38;2;171;159;152m9[0m[38;2;255;242;231m@[0m[38;2;255;237;226m@[0m[38;2;254;236;225m@[0m[38;2;255;237;226m@[0m[38;2;244;227;216m@[0m[38;2;81;76;74m3[0m[38;2;3;4;4m.[0m[38;2;0;0;0m [0m[38;2;74;71;70m5[0m[38;2;183;172;165mB[0m[38;2;243;227;216m@[0m[38;2;255;244;232m@[0m[38;2;255;243;232m@[0m[38;2;255;242;230m@[0m[38;2;255;238;226m@[0m[38;2;255;243;231m@[0m[38;2;188;175;167mB[0m[38;2;19;18;19m;[0m[38;2;185;188;191m&[0m[38;2;245;248;253m@[0m[38;2;241;244;248m@[0m[38;2;240;243;248m@[0m[38;2;247;250;255m@[0m[38;2;173;175;178mB[0m[38;2;22;20;18m;[0m[38;2;154;139;131m#[0m[38;2;208;194;185m&[0m[38;2;23;21;21m;[0m[38;2;165;166;170mB[0m[38;2;247;250;254m@[0m[38;2;143;144;146m#[0m[38;2;11;11;10m,[0m[38;2;87;86;87mh[0m[38;2;198;197;199m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;236;235;240m@[0m[38;2;105;104;111mH[0m[38;2;56;56;59mA[0m[38;2;226;226;229m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;144;144;146m#[0m[38;2;34;31;30mr[0m[38;2;232;216;206m@[0m[38;2;255;238;227m@[0m[38;2;255;239;228m@[0m[38;2;220;205;197m@[0m[38;2;21;20;20m;[0m[38;2;36;34;26mr[0m[38;2;84;79;75m3[0m[38;2;125;117;112mG[0m[38;2;160;149;142m9[0m[38;2;199;185;176m&[0m[38;2;220;205;194m&[0m[38;2;237;220;208m@[0m[38;2;242;226;216m@[0m[38;2;250;232;221m@[0m[38;2;253;235;224m@[0m[38;2;255;239;228m@[0m[38;2;229;212;203m@[0m[38;2;28;27;27mr[0m[38;2;166;153;127mM[0m[38;2;255;254;236m2[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m");
    $display("[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;251;251;251m.[0m[38;2;201;201;201m.[0m[38;2;127;127;127m,[0m[38;2;83;83;84ms[0m[38;2;105;105;108mH[0m[38;2;174;176;180mB[0m[38;2;228;231;236m@[0m[38;2;249;252;255m@[0m[38;2;190;195;205m&[0m[38;2;14;15;19m:[0m[38;2;129;131;135mS[0m[38;2;244;247;252m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;236;239;244m@[0m[38;2;239;242;247m@[0m[38;2;95;98;104mM[0m[38;2;9;9;11m,[0m[38;2;32;32;31mr[0m[38;2;218;198;188m@[0m[38;2;255;232;220m@[0m[38;2;255;229;217m@[0m[38;2;255;229;218m@[0m[38;2;248;218;207m@[0m[38;2;170;155;147m9[0m[38;2;75;70;68m5[0m[38;2;44;40;39ms[0m[38;2;121;112;107mG[0m[38;2;228;213;204m@[0m[38;2;253;237;226m@[0m[38;2;245;227;217m@[0m[38;2;251;233;222m@[0m[38;2;253;235;224m@[0m[38;2;254;236;225m@[0m[38;2;252;234;223m@[0m[38;2;217;199;189m@[0m[38;2;159;142;135m#[0m[38;2;93;80;77mh[0m[38;2;54;45;43mX[0m[38;2;87;77;74m3[0m[38;2;234;205;194m@[0m[38;2;255;220;209m@[0m[38;2;253;219;207m@[0m[38;2;254;223;211m@[0m[38;2;245;221;211m@[0m[38;2;59;56;55mA[0m[38;2;93;94;97mM[0m[38;2;240;243;248m@[0m[38;2;236;239;244m@[0m[38;2;235;238;243m@[0m[38;2;238;241;246m@[0m[38;2;227;230;235m@[0m[38;2;48;50;51mX[0m[38;2;113;86;77mM[0m[38;2;255;246;234m@[0m[38;2;230;215;205m@[0m[38;2;26;25;25m;[0m[38;2;104;104;107mM[0m[38;2;76;76;78m3[0m[38;2;72;72;73m5[0m[38;2;188;188;189m&[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;187;186;189m&[0m[38;2;10;10;11m,[0m[38;2;167;168;172mB[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;243;243;244m@[0m[38;2;42;43;45ms[0m[38;2;131;121;116mS[0m[38;2;255;244;232m@[0m[38;2;253;235;224m@[0m[38;2;255;243;232m@[0m[38;2;157;145;138m9[0m[38;2;41;39;24mr[0m[38;2;188;177;102m9[0m[38;2;26;24;13m;[0m[38;2;11;10;10m,[0m[38;2;71;66;64m2[0m[38;2;142;134;128m#[0m[38;2;190;178;169mB[0m[38;2;220;205;196m@[0m[38;2;237;220;210m@[0m[38;2;250;232;222m@[0m[38;2;255;237;225m@[0m[38;2;255;241;229m@[0m[38;2;176;165;161mB[0m[38;2;83;74;57m2[0m[38;2;249;232;193mS[0m[38;2;255;252;244mr[0m[38;2;255;255;255m.[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m");
    $display("[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m.[0m[38;2;219;219;219m.[0m[38;2;144;144;144m,[0m[38;2;84;83;84mr[0m[38;2;92;92;94mh[0m[38;2;154;156;159mB[0m[38;2;215;217;222m@[0m[38;2;242;245;250m@[0m[38;2;241;245;250m@[0m[38;2;240;242;247m@[0m[38;2;214;219;229m@[0m[38;2;100;109;126mG[0m[38;2;10;10;11m,[0m[38;2;186;189;194m&[0m[38;2;241;244;249m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;240;242;247m@[0m[38;2;202;206;212m@[0m[38;2;23;24;27mi[0m[38;2;49;54;63mA[0m[38;2;0;1;3m.[0m[38;2;83;70;68m5[0m[38;2;255;205;193m@[0m[38;2;255;201;190m@[0m[38;2;252;199;189m@[0m[38;2;165;131;123m#[0m[38;2;116;91;85mM[0m[38;2;172;140;132m9[0m[38;2;239;207;197m@[0m[38;2;255;237;225m@[0m[38;2;255;240;229m@[0m[38;2;250;232;222m@[0m[38;2;157;147;143m9[0m[38;2;241;224;214m@[0m[38;2;255;244;232m@[0m[38;2;255;239;228m@[0m[38;2;251;232;219m@[0m[38;2;255;225;213m@[0m[38;2;255;223;211m@[0m[38;2;255;210;199m@[0m[38;2;248;196;185m@[0m[38;2;238;183;174m&[0m[38;2;232;148;147mB[0m[38;2;252;192;182m@[0m[38;2;255;202;191m@[0m[38;2;255;213;201m@[0m[38;2;135;113;108mG[0m[38;2;32;34;35mr[0m[38;2;212;214;219m@[0m[38;2;239;242;247m@[0m[38;2;235;238;243m@[0m[38;2;237;240;245m@[0m[38;2;241;245;249m@[0m[38;2;108;110;113mH[0m[38;2;51;37;32ms[0m[38;2;208;158;150mB[0m[38;2;167;157;151m9[0m[38;2;76;71;69m5[0m[38;2;4;4;5m.[0m[38;2;47;46;47mX[0m[38;2;163;163;164mB[0m[38;2;251;251;252m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;92;92;94mM[0m[38;2;67;67;68m2[0m[38;2;252;252;252m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;167;167;169mB[0m[38;2;19;18;18m:[0m[38;2;214;200;191m@[0m[38;2;255;240;229m@[0m[38;2;254;239;227m@[0m[38;2;244;209;199m@[0m[38;2;52;39;37ms[0m[38;2;78;74;44m2[0m[38;2;108;101;60mh[0m[38;2;7;6;5m,[0m[38;2;112;104;97mH[0m[38;2;196;182;176m&[0m[38;2;226;210;203m@[0m[38;2;238;222;214m@[0m[38;2;241;224;216m@[0m[38;2;243;226;217m@[0m[38;2;246;229;218m@[0m[38;2;246;231;221m@[0m[38;2;203;190;182m&[0m[38;2;47;44;40mX[0m[38;2;214;190;140m9[0m[38;2;255;246;215mM[0m[38;2;255;253;250m:[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m");
    $display("[38;2;234;234;234m5[0m[38;2;233;233;233m5[0m[38;2;246;246;246m3[0m[38;2;255;255;255m,[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;253;253;253ms[0m[38;2;240;239;239m5[0m[38;2;244;244;244m5[0m[38;2;243;243;242mA[0m[38;2;181;181;180m,[0m[38;2;99;99;100m;[0m[38;2;78;78;79m5[0m[38;2;132;134;136m#[0m[38;2;202;205;209m@[0m[38;2;239;242;247m@[0m[38;2;243;246;251m@[0m[38;2;238;241;246m@[0m[38;2;235;238;243m@[0m[38;2;237;240;244m@[0m[38;2;224;227;234m@[0m[38;2;143;157;181m9[0m[38;2;62;69;82m5[0m[38;2;30;31;34mr[0m[38;2;219;222;229m@[0m[38;2;238;241;246m@[0m[38;2;235;238;243m@[0m[38;2;236;239;244m@[0m[38;2;235;238;243m@[0m[38;2;86;87;89mh[0m[38;2;15;14;15m:[0m[38;2;112;103;99mH[0m[38;2;113;102;97mH[0m[38;2;174;143;136m9[0m[38;2;254;208;197m@[0m[38;2;254;206;195m@[0m[38;2;254;206;195m@[0m[38;2;255;209;197m@[0m[38;2;255;217;206m@[0m[38;2;255;222;211m@[0m[38;2;255;225;213m@[0m[38;2;253;232;220m@[0m[38;2;235;218;208m@[0m[38;2;189;176;169mB[0m[38;2;161;148;140m9[0m[38;2;151;134;129m#[0m[38;2;143;125;119mS[0m[38;2;137;111;109mG[0m[38;2;133;101;98mH[0m[38;2;105;80;76mh[0m[38;2;159;138;132m#[0m[38;2;255;214;203m@[0m[38;2;255;211;200m@[0m[38;2;250;195;186m@[0m[38;2;218;116;121m9[0m[38;2;245;185;178m@[0m[38;2;255;221;209m@[0m[38;2;186;158;151mB[0m[38;2;22;20;20m;[0m[38;2;167;169;173mB[0m[38;2;242;246;251m@[0m[38;2;235;238;243m@[0m[38;2;237;240;245m@[0m[38;2;234;237;242m@[0m[38;2;130;131;135mS[0m[38;2;2;2;2m.[0m[38;2;47;40;38ms[0m[38;2;53;46;48mX[0m[38;2;51;51;55mA[0m[38;2;112;113;117mH[0m[38;2;162;162;164m9[0m[38;2;238;238;239m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;225;226;226m@[0m[38;2;24;24;25m;[0m[38;2;167;167;168mB[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;209;209;212m@[0m[38;2;29;30;32mi[0m[38;2;52;45;42mX[0m[38;2;255;229;218m@[0m[38;2;255;243;232m@[0m[38;2;255;230;220m@[0m[38;2;156;118;109mS[0m[38;2;0;0;0m [0m[38;2;76;71;44m2[0m[38;2;153;143;84mS[0m[38;2;78;73;45m2[0m[38;2;70;67;40m2[0m[38;2;45;43;27ms[0m[38;2;56;53;38mX[0m[38;2;81;77;57m5[0m[38;2;87;82;63m3[0m[38;2;79;75;60m5[0m[38;2;56;53;51mA[0m[38;2;115;108;105mH[0m[38;2;144;135;130m#[0m[38;2;127;113;82mH[0m[38;2;254;229;175mB[0m[38;2;255;247;229m2[0m[38;2;255;255;254m.[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m");
    $display("[38;2;214;214;215mG[0m[38;2;213;212;213mG[0m[38;2;241;241;241mS[0m[38;2;255;255;255m,[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m5[0m[38;2;211;210;210mS[0m[38;2;119;118;118mM[0m[38;2;69;69;68m2[0m[38;2;92;93;95mM[0m[38;2;171;173;177m&[0m[38;2;231;234;239m@[0m[38;2;244;247;252m@[0m[38;2;238;241;246m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;239;241;245m@[0m[38;2;177;185;200m&[0m[38;2;123;140;167m#[0m[38;2;39;42;50ms[0m[38;2;74;75;79m3[0m[38;2;239;242;248m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;236;239;244m@[0m[38;2;236;239;244m@[0m[38;2;67;67;70m5[0m[38;2;7;6;6m,[0m[38;2;120;109;104mH[0m[38;2;228;208;197m@[0m[38;2;255;240;227m@[0m[38;2;255;237;225m@[0m[38;2;255;233;221m@[0m[38;2;254;231;219m@[0m[38;2;253;230;219m@[0m[38;2;253;231;219m@[0m[38;2;252;232;221m@[0m[38;2;253;234;223m@[0m[38;2;255;243;231m@[0m[38;2;136;129;124mS[0m[38;2;83;47;47m2[0m[38;2;202;106;111m#[0m[38;2;205;106;112m#[0m[38;2;214;120;123m9[0m[38;2;227;136;138mB[0m[38;2;242;158;157m&[0m[38;2;154;102;101mG[0m[38;2;78;74;71m5[0m[38;2;255;234;223m@[0m[38;2;253;230;219m@[0m[38;2;252;230;219m@[0m[38;2;253;230;219m@[0m[38;2;255;241;229m@[0m[38;2;214;196;187m&[0m[38;2;34;32;32mr[0m[38;2;130;131;135mS[0m[38;2;242;245;251m@[0m[38;2;235;238;243m@[0m[38;2;237;240;245m@[0m[38;2;242;245;250m@[0m[38;2;97;98;100mM[0m[38;2;15;15;16m:[0m[38;2;114;112;121mG[0m[38;2;157;154;169m9[0m[38;2;179;177;190m&[0m[38;2;225;224;230m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;153;152;154m9[0m[38;2;33;33;34mr[0m[38;2;237;237;238m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;142;142;146m#[0m[38;2;0;0;0m [0m[38;2;29;22;18m;[0m[38;2;190;144;134m9[0m[38;2;175;143;133m9[0m[38;2;130;99;93mH[0m[38;2;36;27;27mi[0m[38;2;7;7;4m,[0m[38;2;143;135;80mG[0m[38;2;215;207;118m&[0m[38;2;254;244;138m@[0m[38;2;255;246;139m@[0m[38;2;244;233;132m@[0m[38;2;244;232;131m@[0m[38;2;248;236;133m@[0m[38;2;247;242;136m@[0m[38;2;170;162;90m#[0m[38;2;18;16;15m:[0m[38;2;82;78;76m3[0m[38;2;81;73;54m5[0m[38;2;210;184;125mB[0m[38;2;255;238;196mS[0m[38;2;255;251;243mi[0m[38;2;255;255;255m:[0m[38;2;243;243;243mh[0m[38;2;229;229;229m3[0m[38;2;232;232;232m5[0m[38;2;235;235;235m5[0m[38;2;237;237;237m5[0m[38;2;238;238;239m2[0m[38;2;240;240;241m2[0m[38;2;242;242;241m2[0m");
    $display("[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;247;247;247m.[0m[38;2;159;159;158m,[0m[38;2;70;70;70mi[0m[38;2;104;105;107mH[0m[38;2;195;197;202m&[0m[38;2;241;244;249m@[0m[38;2;243;246;251m@[0m[38;2;229;231;237m@[0m[38;2;222;224;230m@[0m[38;2;232;235;240m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;237;240;244m@[0m[38;2;224;227;234m@[0m[38;2;136;150;174m9[0m[38;2;121;137;163m#[0m[38;2;23;26;30mi[0m[38;2;116;116;118mG[0m[38;2;244;246;251m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;240;243;248m@[0m[38;2;194;196;200m&[0m[38;2;22;22;23m;[0m[38;2;76;84;99mh[0m[38;2;48;55;65mA[0m[38;2;34;34;37mr[0m[38;2;86;81;78m3[0m[38;2;162;152;145m9[0m[38;2;219;204;195m@[0m[38;2;250;233;223m@[0m[38;2;255;243;232m@[0m[38;2;255;244;233m@[0m[38;2;255;242;230m@[0m[38;2;255;239;228m@[0m[38;2;255;241;230m@[0m[38;2;206;193;184m&[0m[38;2;72;54;52mA[0m[38;2;192;105;109m#[0m[38;2;252;169;167m&[0m[38;2;255;182;177m@[0m[38;2;255;185;180m@[0m[38;2;255;190;185m@[0m[38;2;120;90;88mM[0m[38;2;131;125;120mS[0m[38;2;255;244;233m@[0m[38;2;255;238;227m@[0m[38;2;255;241;229m@[0m[38;2;255;243;232m@[0m[38;2;193;182;174m&[0m[38;2;37;34;34mr[0m[38;2;107;108;112mH[0m[38;2;239;242;247m@[0m[38;2;236;239;244m@[0m[38;2;238;241;246m@[0m[38;2;240;243;248m@[0m[38;2;126;127;130mS[0m[38;2;27;27;29mi[0m[38;2;142;140;151m#[0m[38;2;197;194;210m&[0m[38;2;216;214;224m@[0m[38;2;245;245;247m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;144;144;145m#[0m[38;2;39;39;40ms[0m[38;2;229;229;230m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;253;253;254m@[0m[38;2;252;252;254m@[0m[38;2;253;253;255m@[0m[38;2;241;241;245m@[0m[38;2;183;181;195m&[0m[38;2;125;123;132mS[0m[38;2;74;74;79m3[0m[38;2;22;22;22m;[0m[38;2;6;5;3m.[0m[38;2;2;3;0m.[0m[38;2;113;108;63mM[0m[38;2;209;201;115mB[0m[38;2;254;243;138m@[0m[38;2;255;249;141m@[0m[38;2;255;247;140m@[0m[38;2;255;244;139m@[0m[38;2;255;245;139m@[0m[38;2;255;245;139m@[0m[38;2;255;244;139m@[0m[38;2;255;253;143m@[0m[38;2;162;154;89m#[0m[38;2;0;0;1m.[0m[38;2;136;119;77mH[0m[38;2;244;213;140m@[0m[38;2;255;227;162m&[0m[38;2;255;241;214mh[0m[38;2;255;254;252m,[0m[38;2;255;255;255m;[0m[38;2;237;237;237mS[0m[38;2;213;212;213mG[0m[38;2;213;213;214mG[0m[38;2;214;214;214mG[0m[38;2;213;213;213mS[0m[38;2;212;212;213mS[0m[38;2;213;213;214mS[0m[38;2;218;218;217m#[0m");
    $display("[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m.[0m[38;2;190;190;190m:[0m[38;2;69;69;69m;[0m[38;2;87;88;90mM[0m[38;2;195;198;202m@[0m[38;2;242;245;250m@[0m[38;2;242;245;249m@[0m[38;2;235;238;243m@[0m[38;2;207;212;221m@[0m[38;2;215;218;225m@[0m[38;2;234;237;242m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;239;242;246m@[0m[38;2;184;192;206m&[0m[38;2;125;142;170m#[0m[38;2;106;119;141mS[0m[38;2;7;8;9m,[0m[38;2;144;145;149m#[0m[38;2;243;246;251m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;243;246;251m@[0m[38;2;128;128;131mS[0m[38;2;20;22;26m;[0m[38;2;123;139;164m#[0m[38;2;129;146;173m9[0m[38;2;116;131;155m#[0m[38;2;68;77;92m3[0m[38;2;2;2;3m.[0m[38;2;19;19;20m;[0m[38;2;54;52;51mA[0m[38;2;100;94;90mM[0m[38;2;149;139;133m#[0m[38;2;190;177;169m&[0m[38;2;224;209;199m@[0m[38;2;243;226;215m@[0m[38;2;255;240;229m@[0m[38;2;218;205;196m@[0m[38;2;158;138;129m#[0m[38;2;246;189;182m@[0m[38;2;255;198;192m@[0m[38;2;255;199;192m@[0m[38;2;255;206;199m@[0m[38;2;216;187;179m&[0m[38;2;235;219;209m@[0m[38;2;244;228;217m@[0m[38;2;234;218;208m@[0m[38;2;218;205;197m@[0m[38;2;136;127;121mS[0m[38;2;8;8;7m,[0m[38;2;98;100;103mM[0m[38;2;235;238;243m@[0m[38;2;237;240;245m@[0m[38;2;240;243;248m@[0m[38;2;230;233;239m@[0m[38;2;101;102;105mH[0m[38;2;34;33;36mr[0m[38;2;158;155;166m9[0m[38;2;218;216;225m@[0m[38;2;241;241;243m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;243;244;244m@[0m[38;2;128;128;130mS[0m[38;2;66;66;68m2[0m[38;2;108;108;110mH[0m[38;2;146;145;151m9[0m[38;2;170;168;178mB[0m[38;2;153;151;163m9[0m[38;2;125;125;135mS[0m[38;2;102;101;107mH[0m[38;2;104;100;98mM[0m[38;2;83;81;79m3[0m[38;2;35;35;41mr[0m[38;2;34;32;27mi[0m[38;2;86;81;48m5[0m[38;2;205;196;112mB[0m[38;2;255;255;146m@[0m[38;2;255;255;146m@[0m[38;2;255;251;142m@[0m[38;2;249;237;134m@[0m[38;2;238;226;129m&[0m[38;2;255;246;140m@[0m[38;2;255;246;139m@[0m[38;2;255;243;138m@[0m[38;2;255;243;138m@[0m[38;2;255;252;143m@[0m[38;2;161;152;87mS[0m[38;2;0;0;2m.[0m[38;2;209;181;120mB[0m[38;2;255;225;150m@[0m[38;2;254;228;176m9[0m[38;2;255;248;235mX[0m[38;2;255;255;255m.[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m");
    $display("[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;245;245;245m,[0m[38;2;116;116;116m:[0m[38;2;51;52;53mA[0m[38;2;165;166;170mB[0m[38;2;240;243;248m@[0m[38;2;240;243;249m@[0m[38;2;238;241;245m@[0m[38;2;228;231;237m@[0m[38;2;181;188;202m&[0m[38;2;210;214;222m@[0m[38;2;237;240;245m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;236;239;244m@[0m[38;2;231;233;239m@[0m[38;2;145;159;182mB[0m[38;2;107;120;143mS[0m[38;2;34;36;41mr[0m[38;2;7;7;7m,[0m[38;2;153;154;159m9[0m[38;2;244;247;252m@[0m[38;2;236;239;244m@[0m[38;2;235;238;243m@[0m[38;2;242;245;250m@[0m[38;2;85;85;87mh[0m[38;2;42;46;54mX[0m[38;2;129;145;172m9[0m[38;2;127;144;170m9[0m[38;2;113;127;150mS[0m[38;2;56;62;73m2[0m[38;2;3;3;3m.[0m[38;2;32;34;37mr[0m[38;2;32;32;35mr[0m[38;2;28;28;31mi[0m[38;2;36;36;39mr[0m[38;2;51;51;54mA[0m[38;2;27;26;26mi[0m[38;2;60;58;58mA[0m[38;2;93;88;87mh[0m[38;2;119;111;109mG[0m[38;2;125;117;113mG[0m[38;2;111;102;98mH[0m[38;2;111;101;97mH[0m[38;2;112;103;99mH[0m[38;2;106;100;96mM[0m[38;2;97;92;89mM[0m[38;2;81;77;75m3[0m[38;2;73;70;69m5[0m[38;2;40;39;39ms[0m[38;2;9;8;8m,[0m[38;2;0;0;0m [0m[38;2;117;118;121mG[0m[38;2;238;241;246m@[0m[38;2;238;241;246m@[0m[38;2;243;246;251m@[0m[38;2;210;212;217m@[0m[38;2;67;67;69m5[0m[38;2;60;59;62m2[0m[38;2;195;194;200m&[0m[38;2;247;246;249m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;251;251;252m@[0m[38;2;252;253;253m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;225;225;226m@[0m[38;2;144;143;149m#[0m[38;2;89;88;95mh[0m[38;2;14;15;17m:[0m[38;2;61;55;44mA[0m[38;2;154;135;91mS[0m[38;2;184;161;106m9[0m[38;2;125;108;69mM[0m[38;2;33;30;17mi[0m[38;2;114;107;62mM[0m[38;2;228;219;125m&[0m[38;2;255;250;142m@[0m[38;2;235;224;128m&[0m[38;2;189;180;103m9[0m[38;2;145;137;80mG[0m[38;2;100;95;56mh[0m[38;2;78;73;47m2[0m[38;2;42;39;26mr[0m[38;2;106;100;58mh[0m[38;2;241;232;132m@[0m[38;2;255;245;139m@[0m[38;2;255;243;138m@[0m[38;2;255;250;142m@[0m[38;2;182;173;100m9[0m[38;2;14;13;11m:[0m[38;2;207;180;117mB[0m[38;2;255;225;154m@[0m[38;2;254;236;198mG[0m[38;2;255;253;249m;[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m");
    $display("[38;2;255;255;255m [0m[38;2;233;233;233m,[0m[38;2;73;73;73m:[0m[38;2;77;77;80mh[0m[38;2;217;219;224m@[0m[38;2;243;246;251m@[0m[38;2;236;239;244m@[0m[38;2;239;241;246m@[0m[38;2;216;220;228m@[0m[38;2;155;165;184mB[0m[38;2;203;208;218m@[0m[38;2;239;241;246m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;238;241;246m@[0m[38;2;202;208;219m@[0m[38;2;120;136;161m#[0m[38;2;33;35;41mr[0m[38;2;57;61;69m2[0m[38;2;32;32;34mr[0m[38;2;139;140;143m#[0m[38;2;245;248;253m@[0m[38;2;230;233;238m@[0m[38;2;236;239;244m@[0m[38;2;239;242;247m@[0m[38;2;70;70;72m5[0m[38;2;53;58;68m2[0m[38;2;131;148;175m9[0m[38;2;113;126;149mS[0m[38;2;26;28;31mi[0m[38;2;95;94;98mM[0m[38;2;32;32;34mr[0m[38;2;49;49;50mX[0m[38;2;166;164;176mB[0m[38;2;168;165;179mB[0m[38;2;159;156;169m9[0m[38;2;135;133;140m#[0m[38;2;2;2;2m.[0m[38;2;79;78;83m3[0m[38;2;164;161;175mB[0m[38;2;139;137;148m#[0m[38;2;28;29;31mi[0m[38;2;28;29;30mi[0m[38;2;99;98;105mM[0m[38;2;35;36;38mr[0m[38;2;31;32;33mr[0m[38;2;119;118;128mG[0m[38;2;157;154;168m9[0m[38;2;112;110;118mG[0m[38;2;8;8;9m,[0m[38;2;12;11;12m,[0m[38;2;142;144;147m#[0m[38;2;241;243;248m@[0m[38;2;239;243;248m@[0m[38;2;242;244;250m@[0m[38;2;168;169;172mB[0m[38;2;34;34;35mr[0m[38;2;110;109;111mH[0m[38;2;238;238;239m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;240;240;242m@[0m[38;2;211;211;218m@[0m[38;2;207;205;214m@[0m[38;2;215;213;223m@[0m[38;2;220;218;227m@[0m[38;2;219;218;226m@[0m[38;2;223;223;228m@[0m[38;2;232;231;234m@[0m[38;2;239;239;241m@[0m[38;2;248;249;250m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;105;105;110mH[0m[38;2;46;42;37mr[0m[38;2;235;210;154mB[0m[38;2;234;207;139m&[0m[38;2;84;74;49m5[0m[38;2;46;43;26ms[0m[38;2;145;137;80mG[0m[38;2;182;174;101m9[0m[38;2;143;137;80mG[0m[38;2;100;95;56mh[0m[38;2;71;67;40m2[0m[38;2;86;82;48m5[0m[38;2;120;114;67mM[0m[38;2;163;155;89m#[0m[38;2;211;204;118mB[0m[38;2;175;166;97m#[0m[38;2;2;2;3m.[0m[38;2;150;141;83mS[0m[38;2;255;252;143m@[0m[38;2;255;243;138m@[0m[38;2;255;251;142m@[0m[38;2;175;167;96m#[0m[38;2;26;23;17m;[0m[38;2;227;197;131m&[0m[38;2;255;229;170mB[0m[38;2;255;245;226m2[0m[38;2;255;255;255m.[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m");
    $display("[38;2;242;242;242m,[0m[38;2;71;71;71m:[0m[38;2;80;80;82mh[0m[38;2;233;236;240m@[0m[38;2;240;243;248m@[0m[38;2;235;238;243m@[0m[38;2;239;241;246m@[0m[38;2;201;206;216m@[0m[38;2;133;147;171m9[0m[38;2;180;188;202m&[0m[38;2;239;242;246m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;238;240;244m@[0m[38;2;168;178;197m&[0m[38;2;70;79;93m3[0m[38;2;21;22;24m;[0m[38;2;121;136;160m#[0m[38;2;51;54;62mA[0m[38;2;105;105;106mH[0m[38;2;119;120;122mG[0m[38;2;120;121;124mG[0m[38;2;241;245;250m@[0m[38;2;242;245;250m@[0m[38;2;72;73;75m5[0m[38;2;52;58;69m2[0m[38;2;133;150;177m9[0m[38;2;53;59;69m2[0m[38;2;36;35;36mr[0m[38;2;129;130;132mS[0m[38;2;18;18;19m:[0m[38;2;48;46;45mX[0m[38;2;95;92;92mM[0m[38;2;103;99;98mM[0m[38;2;71;67;65m5[0m[38;2;11;11;11m,[0m[38;2;14;14;14m:[0m[38;2;23;23;24m;[0m[38;2;66;66;69m5[0m[38;2;23;23;24m;[0m[38;2;38;38;38ms[0m[38;2;21;21;21m;[0m[38;2;26;26;28mi[0m[38;2;95;95;100mM[0m[38;2;15;15;16m:[0m[38;2;20;20;20m;[0m[38;2;39;38;41ms[0m[38;2;37;41;48ms[0m[38;2;112;117;129mG[0m[38;2;186;188;192m&[0m[38;2;242;245;250m@[0m[38;2;242;245;250m@[0m[38;2;228;231;236m@[0m[38;2;111;111;114mG[0m[38;2;30;30;31mi[0m[38;2;18;18;19m:[0m[38;2;127;126;128mS[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;246;246;249m@[0m[38;2;223;221;229m@[0m[38;2;196;193;207m&[0m[38;2;171;167;182mB[0m[38;2;143;140;153m9[0m[38;2;111;109;119mG[0m[38;2;82;81;87m3[0m[38;2;82;82;85m2[0m[38;2;127;127;130mA[0m[38;2;144;144;148m5[0m[38;2;117;117;120mM[0m[38;2;110;109;110mH[0m[38;2;113;112;111mH[0m[38;2;126;126;128mS[0m[38;2;142;142;142m9[0m[38;2;114;114;115mG[0m[38;2;45;43;41mi[0m[38;2;211;192;155mS[0m[38;2;189;171;121m#[0m[38;2;45;40;27mr[0m[38;2;18;18;12m:[0m[38;2;90;85;51m3[0m[38;2;118;112;67mM[0m[38;2;142;135;79mG[0m[38;2;187;178;103m9[0m[38;2;226;215;123m&[0m[38;2;253;241;137m@[0m[38;2;255;255;145m@[0m[38;2;255;255;146m@[0m[38;2;255;255;145m@[0m[38;2;255;253;144m@[0m[38;2;255;255;145m@[0m[38;2;76;72;44m2[0m[38;2;89;84;51m5[0m[38;2;255;249;142m@[0m[38;2;255;243;138m@[0m[38;2;255;251;142m@[0m[38;2;136;128;75mG[0m[38;2;42;37;26mr[0m[38;2;243;210;142m&[0m[38;2;254;233;190m9[0m[38;2;255;252;245mX[0m[38;2;255;255;255m,[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m");
    $display("[38;2;131;131;131m;[0m[38;2;36;36;37mX[0m[38;2;218;220;225m@[0m[38;2;240;243;248m@[0m[38;2;236;239;243m@[0m[38;2;238;240;245m@[0m[38;2;191;197;210m&[0m[38;2;124;140;166m#[0m[38;2;148;160;181mB[0m[38;2;232;234;240m@[0m[38;2;236;239;244m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;236;239;244m@[0m[38;2;228;231;237m@[0m[38;2;130;142;163m#[0m[38;2;20;21;24m;[0m[38;2;72;79;93m3[0m[38;2;133;150;178m9[0m[38;2;94;105;124mH[0m[38;2;38;40;44ms[0m[38;2;5;5;6m.[0m[38;2;84;84;87mh[0m[38;2;242;245;251m@[0m[38;2;249;252;255m@[0m[38;2;102;103;105mH[0m[38;2;26;29;35mi[0m[38;2;99;110;129mG[0m[38;2;24;24;25m;[0m[38;2;69;69;70m5[0m[38;2;123;114;110mG[0m[38;2;204;190;182m&[0m[38;2;230;214;203m@[0m[38;2;241;224;213m@[0m[38;2;255;240;228m@[0m[38;2;172;160;153mB[0m[38;2;66;63;61m2[0m[38;2;67;65;64m2[0m[38;2;7;7;7m,[0m[38;2;25;25;26mi[0m[38;2;58;57;59mA[0m[38;2;43;43;44ms[0m[38;2;34;34;36mr[0m[38;2;28;28;30mi[0m[38;2;114;112;119mG[0m[38;2;25;24;25m;[0m[38;2;33;37;44ms[0m[38;2;83;93;112mM[0m[38;2;167;177;192m&[0m[38;2;237;240;246m@[0m[38;2;243;246;251m@[0m[38;2;245;248;253m@[0m[38;2;197;199;203m&[0m[38;2;67;67;69m5[0m[38;2;24;24;27mi[0m[38;2;46;46;51mX[0m[38;2;17;17;17m:[0m[38;2;95;95;97mM[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;238;238;241m@[0m[38;2;197;195;203m&[0m[38;2;151;148;159m9[0m[38;2;100;98;107mH[0m[38;2;70;69;73m3[0m[38;2;83;83;84m2[0m[38;2;115;114;113mi[0m[38;2;153;153;154mh[0m[38;2;166;166;166mB[0m[38;2;178;178;178m#[0m[38;2;242;242;242mH[0m[38;2;255;255;255mi[0m[38;2;245;245;245m.[0m[38;2;231;231;230m:[0m[38;2;217;216;214m,[0m[38;2;200;200;200m.[0m[38;2;185;185;185m.[0m[38;2;178;176;173ms[0m[38;2;221;206;181m9[0m[38;2;254;228;170m&[0m[38;2;107;92;65mh[0m[38;2;20;19;13m;[0m[38;2;162;154;89m#[0m[38;2;247;238;135m@[0m[38;2;255;255;146m@[0m[38;2;255;244;139m@[0m[38;2;186;177;102m9[0m[38;2;161;152;88m#[0m[38;2;148;140;82mS[0m[38;2;134;126;74mG[0m[38;2;123;116;68mH[0m[38;2;115;109;66mM[0m[38;2;91;87;53m3[0m[38;2;136;130;76mG[0m[38;2;142;134;79mG[0m[38;2;36;34;23mr[0m[38;2;238;227;129m&[0m[38;2;255;246;140m@[0m[38;2;255;248;140m@[0m[38;2;81;77;46m5[0m[38;2;87;75;51m5[0m[38;2;252;222;154m@[0m[38;2;227;210;183m&[0m[38;2;208;207;208mB[0m[38;2;210;210;211m9[0m[38;2;217;217;217m#[0m[38;2;224;223;224mG[0m[38;2;233;233;233mM[0m[38;2;241;241;241m5[0m[38;2;247;247;247mA[0m[38;2;252;252;252mr[0m[38;2;253;253;253m:[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m");
    $display("[38;2;32;32;32m:[0m[38;2;119;120;123mS[0m[38;2;244;247;252m@[0m[38;2;236;239;244m@[0m[38;2;237;240;244m@[0m[38;2;185;192;206m&[0m[38;2;126;142;168m#[0m[38;2;126;141;167m#[0m[38;2;209;214;223m@[0m[38;2;238;241;246m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;238;241;245m@[0m[38;2;209;215;226m@[0m[38;2;83;91;107mM[0m[38;2;15;15;17m:[0m[38;2;113;127;149mS[0m[38;2;127;143;170m9[0m[38;2;126;143;169m#[0m[38;2;113;127;151mS[0m[38;2;96;108;128mH[0m[38;2;58;63;72m2[0m[38;2;92;94;98mM[0m[38;2;185;186;189m&[0m[38;2;159;162;170mB[0m[38;2;18;20;23m;[0m[38;2;38;41;47ms[0m[38;2;126;125;130mS[0m[38;2;183;183;189m&[0m[38;2;38;36;36mr[0m[38;2;149;140;134m#[0m[38;2;255;241;230m@[0m[38;2;255;242;230m@[0m[38;2;254;235;224m@[0m[38;2;255;237;226m@[0m[38;2;254;240;229m@[0m[38;2;196;182;175m&[0m[38;2;4;4;5m.[0m[38;2;5;5;5m.[0m[38;2;25;25;26m;[0m[38;2;17;17;18m:[0m[38;2;44;44;46mX[0m[38;2;5;5;5m.[0m[38;2;35;38;44ms[0m[38;2;89;101;121mH[0m[38;2;132;147;171m9[0m[38;2;194;202;216m@[0m[38;2;244;246;251m@[0m[38;2;246;249;254m@[0m[38;2;230;233;238m@[0m[38;2;142;143;146m#[0m[38;2;24;25;25m;[0m[38;2;0;0;0m [0m[38;2;8;8;9m,[0m[38;2;76;75;80m3[0m[38;2;122;121;131mS[0m[38;2;222;222;227m@[0m[38;2;244;244;245m@[0m[38;2;192;192;194m&[0m[38;2;125;125;129mS[0m[38;2;79;78;82m3[0m[38;2;50;49;52mA[0m[38;2;21;21;22m;[0m[38;2;95;94;93ms[0m[38;2;176;176;177mS[0m[38;2;251;250;249m#[0m[38;2;255;255;255mi[0m[38;2;255;255;255mr[0m[38;2;248;248;248mG[0m[38;2;203;202;203mB[0m[38;2;175;175;176m&[0m[38;2;194;195;195m&[0m[38;2;237;237;237mS[0m[38;2;255;255;255ms[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255mi[0m[38;2;249;243;233mS[0m[38;2;248;230;192m9[0m[38;2;247;222;169mB[0m[38;2;168;148;107mS[0m[38;2;86;77;50m5[0m[38;2;93;88;51m3[0m[38;2;165;160;91m#[0m[38;2;213;204;117mB[0m[38;2;109;104;61mh[0m[38;2;30;28;20mi[0m[38;2;88;82;51m5[0m[38;2;176;167;97m9[0m[38;2;217;211;120m&[0m[38;2;197;187;108mB[0m[38;2;27;25;18m;[0m[38;2;167;158;92m#[0m[38;2;237;226;130m&[0m[38;2;33;30;21mi[0m[38;2;157;148;87mS[0m[38;2;255;255;145m@[0m[38;2;239;227;130m&[0m[38;2;35;32;21mi[0m[38;2;145;127;88mG[0m[38;2;255;238;187m9[0m[38;2;255;247;234m5[0m[38;2;250;250;250mX[0m[38;2;242;242;242m2[0m[38;2;235;235;235mh[0m[38;2;227;227;227mG[0m[38;2;218;218;219m#[0m[38;2;214;213;214m9[0m[38;2;205;205;206mB[0m[38;2;212;212;213mB[0m[38;2;251;251;250mM[0m[38;2;255;255;255m [0m[38;2;254;254;254m:[0m[38;2;242;242;243mM[0m");
    $display("[38;2;13;13;13m,[0m[38;2;154;156;159m9[0m[38;2;243;246;251m@[0m[38;2;238;241;245m@[0m[38;2;186;194;208m&[0m[38;2;125;141;168m#[0m[38;2;89;101;120mH[0m[38;2;164;173;189mB[0m[38;2;238;240;245m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;239;242;246m@[0m[38;2;183;190;205m&[0m[38;2;41;45;53mX[0m[38;2;43;48;55mX[0m[38;2;127;143;170m9[0m[38;2;125;141;167m#[0m[38;2;125;141;167m#[0m[38;2;127;143;169m9[0m[38;2;128;145;172m9[0m[38;2;126;142;168m#[0m[38;2;103;117;140mG[0m[38;2;86;95;110mM[0m[38;2;95;100;111mH[0m[38;2;61;64;71mA[0m[38;2;61;60;64m2[0m[38;2;103;102;109mH[0m[38;2;51;50;53mX[0m[38;2;100;100;101mM[0m[38;2;63;63;64m2[0m[38;2;94;88;85mh[0m[38;2;221;207;198m@[0m[38;2;255;242;230m@[0m[38;2;255;241;230m@[0m[38;2;255;242;231m@[0m[38;2;245;230;220m@[0m[38;2;103;97;94mM[0m[38;2;6;6;7m,[0m[38;2;52;51;54mA[0m[38;2;66;64;67m2[0m[38;2;24;24;24m;[0m[38;2;17;18;21m;[0m[38;2;87;96;112mM[0m[38;2;171;183;203m&[0m[38;2;226;230;238m@[0m[38;2;240;242;246m@[0m[38;2;182;184;187m&[0m[38;2;115;116;118mG[0m[38;2;55;55;59mA[0m[38;2;18;19;25m;[0m[38;2;1;1;2m.[0m[38;2;1;1;1m.[0m[38;2;8;8;8m,[0m[38;2;79;78;84m3[0m[38;2;193;190;205m&[0m[38;2;146;144;152m9[0m[38;2;78;78;80m3[0m[38;2;91;91;93mh[0m[38;2;78;78;80m3[0m[38;2;53;53;54mA[0m[38;2;73;72;72mr[0m[38;2;150;150;149mX[0m[38;2;209;208;207m;[0m[38;2;181;181;181m;[0m[38;2;156;155;154m3[0m[38;2;148;148;149m#[0m[38;2;246;245;245mS[0m[38;2;255;255;255m [0m[38;2;255;255;255m:[0m[38;2;252;252;252m3[0m[38;2;224;224;224m#[0m[38;2;199;199;201m&[0m[38;2;199;199;200m&[0m[38;2;226;226;227m#[0m[38;2;252;252;251m5[0m[38;2;255;255;255m,[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;254;252m,[0m[38;2;255;250;237mX[0m[38;2;255;248;216mM[0m[38;2;251;230;181m#[0m[38;2;197;177;133m9[0m[38;2;122;108;80mH[0m[38;2;88;79;53m3[0m[38;2;109;103;60mM[0m[38;2;126;119;69mH[0m[38;2;99;93;55m3[0m[38;2;86;81;48m5[0m[38;2;115;110;65mM[0m[38;2;138;130;76mG[0m[38;2;124;116;70mH[0m[38;2;207;196;113mB[0m[38;2;224;218;124m&[0m[38;2;114;107;64mM[0m[38;2;39;36;24mr[0m[38;2;241;231;132m@[0m[38;2;188;178;102m9[0m[38;2;14;13;12m:[0m[38;2;210;189;145m#[0m[38;2;255;244;212mH[0m[38;2;255;253;249m:[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m.[0m[38;2;255;255;255m:[0m[38;2;253;253;253m;[0m[38;2;254;254;254m:[0m[38;2;255;255;255m [0m[38;2;255;255;255m;[0m[38;2;242;242;242mS[0m");
    $display("[38;2;17;17;17m:[0m[38;2;144;145;148m#[0m[38;2;247;250;255m@[0m[38;2;208;213;223m@[0m[38;2;114;127;150mS[0m[38;2;53;58;68m2[0m[38;2;35;37;42ms[0m[38;2;208;212;220m@[0m[38;2;239;242;247m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;239;241;246m@[0m[38;2;154;164;180mB[0m[38;2;16;17;21m:[0m[38;2;69;75;88m3[0m[38;2;130;146;173m9[0m[38;2;125;141;167m#[0m[38;2;125;141;167m#[0m[38;2;125;141;167m#[0m[38;2;125;141;167m#[0m[38;2;125;141;167m#[0m[38;2;127;143;170m9[0m[38;2;129;146;173m9[0m[38;2;94;106;125mH[0m[38;2;33;35;39mr[0m[38;2;70;69;70m5[0m[38;2;83;83;83m3[0m[38;2;24;23;24m;[0m[38;2;223;222;223m@[0m[38;2;252;252;253m@[0m[38;2;86;86;88mh[0m[38;2;32;28;26mi[0m[38;2;186;162;152mB[0m[38;2;203;182;173m&[0m[38;2;210;195;186m&[0m[38;2;200;186;177m&[0m[38;2;66;62;60m2[0m[38;2;38;38;41ms[0m[38;2;79;78;81m3[0m[38;2;73;72;74m5[0m[38;2;35;36;39mr[0m[38;2;45;50;58mX[0m[38;2;93;97;105mM[0m[38;2;145;146;149m9[0m[38;2;163;164;167mB[0m[38;2;94;95;97mM[0m[38;2;14;14;18m:[0m[38;2;12;13;19m:[0m[38;2;24;25;35mi[0m[38;2;27;27;35mi[0m[38;2;6;6;6m,[0m[38;2;18;18;22m;[0m[38;2;25;26;33mi[0m[38;2;13;13;13m:[0m[38;2;68;68;71m5[0m[38;2;63;62;65m2[0m[38;2;177;179;182mB[0m[38;2;130;131;133mS[0m[38;2;39;38;39ms[0m[38;2;43;43;43mi[0m[38;2;76;76;76mi[0m[38;2;63;63;65ms[0m[38;2;44;45;48mX[0m[38;2;46;46;51mA[0m[38;2;43;43;47mX[0m[38;2;7;7;8m;[0m[38;2;179;178;177mX[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255mr[0m[38;2;241;241;240mH[0m[38;2;209;209;210mB[0m[38;2;196;196;196m&[0m[38;2;214;214;215mB[0m[38;2;244;244;243mH[0m[38;2;254;254;254mi[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m.[0m[38;2;255;253;249m;[0m[38;2;255;253;237mA[0m[38;2;255;250;222mH[0m[38;2;247;228;191m#[0m[38;2;200;182;142m#[0m[38;2;150;132;98mG[0m[38;2;112;100;68mM[0m[38;2;89;81;52m3[0m[38;2;73;68;40m2[0m[38;2;64;61;37mA[0m[38;2;42;40;26mr[0m[38;2;13;13;11m:[0m[38;2;19;18;13m:[0m[38;2;31;29;19mi[0m[38;2;18;16;13m:[0m[38;2;96;89;56m3[0m[38;2;74;69;46m2[0m[38;2;103;94;77m5[0m[38;2;252;232;192mS[0m[38;2;255;247;230m2[0m[38;2;255;254;253m,[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m");
    $display("[38;2;65;65;65m;[0m[38;2;83;83;85mh[0m[38;2;235;238;244m@[0m[38;2;137;148;168m9[0m[38;2;32;35;41mr[0m[38;2;60;60;58m;[0m[38;2;20;21;24m;[0m[38;2;169;174;187mB[0m[38;2;240;242;247m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;236;239;244m@[0m[38;2;235;237;243m@[0m[38;2;126;133;149m#[0m[38;2;3;3;3m.[0m[38;2;71;78;90m3[0m[38;2;129;146;173m9[0m[38;2;125;141;167m#[0m[38;2;125;141;167m#[0m[38;2;125;141;167m#[0m[38;2;125;141;167m#[0m[38;2;125;141;167m#[0m[38;2;126;142;169m#[0m[38;2;117;132;155m#[0m[38;2;22;24;28mi[0m[38;2;128;128;128mS[0m[38;2;248;248;248m@[0m[38;2;255;255;255m@[0m[38;2;130;129;130mS[0m[38;2;48;48;49mX[0m[38;2;180;180;182m&[0m[38;2;245;246;246m@[0m[38;2;178;178;179mB[0m[38;2;159;155;155m9[0m[38;2;142;139;139m#[0m[38;2;121;120;121mG[0m[38;2;72;72;73m5[0m[38;2;0;0;1m.[0m[38;2;72;72;78m5[0m[38;2;72;72;79m5[0m[38;2;66;66;73m5[0m[38;2;66;66;73m5[0m[38;2;58;57;62m2[0m[38;2;53;52;56mA[0m[38;2;52;51;56mA[0m[38;2;50;50;55mA[0m[38;2;32;33;41mr[0m[38;2;30;30;40mr[0m[38;2;38;39;48ms[0m[38;2;54;55;63mA[0m[38;2;65;65;72m5[0m[38;2;14;15;16m:[0m[38;2;23;24;31mi[0m[38;2;9;10;11m,[0m[38;2;22;22;26m;[0m[38;2;13;13;14m:[0m[38;2;36;36;37mr[0m[38;2;43;43;45ms[0m[38;2;10;10;12m,[0m[38;2;39;39;43ms[0m[38;2;62;63;68m2[0m[38;2;69;69;76m3[0m[38;2;77;77;86m3[0m[38;2;83;83;91mh[0m[38;2;85;85;94mh[0m[38;2;79;80;87m3[0m[38;2;8;8;9m:[0m[38;2;150;150;151m;[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;252;252;252m;[0m[38;2;254;254;254mi[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m:[0m[38;2;250;250;250m3[0m[38;2;222;222;222m9[0m[38;2;197;197;198m&[0m[38;2;236;236;236m9[0m[38;2;254;254;253mi[0m[38;2;255;255;255m,[0m[38;2;255;255;255m.[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m.[0m[38;2;255;254;250m:[0m[38;2;255;254;241mX[0m[38;2;255;251;225mh[0m[38;2;255;240;204mS[0m[38;2;238;216;173m#[0m[38;2;207;184;137m#[0m[38;2;174;153;111mS[0m[38;2;147;128;91mG[0m[38;2;148;128;88mS[0m[38;2;188;164;114m9[0m[38;2;213;187;133mB[0m[38;2;219;193;140mB[0m[38;2;217;193;147m#[0m[38;2;230;210;170mS[0m[38;2;255;237;202mG[0m[38;2;255;246;225m5[0m[38;2;255;253;248m;[0m[38;2;255;255;255m.[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m");
    $display("[38;2;189;189;188m;[0m[38;2;31;30;30mi[0m[38;2;134;141;154m9[0m[38;2;78;88;105mM[0m[38;2;79;79;78m:[0m[38;2;168;168;168mi[0m[38;2;15;15;18m;[0m[38;2;122;134;155m#[0m[38;2;218;222;230m@[0m[38;2;239;241;246m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;236;239;244m@[0m[38;2;232;236;243m@[0m[38;2;105;113;128mG[0m[38;2;0;0;0m [0m[38;2;67;73;86m3[0m[38;2;130;146;173m9[0m[38;2;125;141;167m#[0m[38;2;126;142;168m#[0m[38;2;126;143;169m#[0m[38;2;126;142;169m#[0m[38;2;126;142;168m#[0m[38;2;127;144;170m9[0m[38;2;113;126;149mS[0m[38;2;12;12;14m:[0m[38;2;178;177;178mB[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;186;186;187m&[0m[38;2;74;74;75m5[0m[38;2;121;120;123mG[0m[38;2;226;226;229m@[0m[38;2;186;186;189m&[0m[38;2;133;133;135m#[0m[38;2;104;103;105mH[0m[38;2;54;54;55mX[0m[38;2;29;29;31mi[0m[38;2;79;79;87m3[0m[38;2;83;83;92mh[0m[38;2;83;83;92mh[0m[38;2;84;84;92mh[0m[38;2;85;85;93mh[0m[38;2;85;85;93mh[0m[38;2;71;71;78m5[0m[38;2;44;45;52mX[0m[38;2;48;49;57mX[0m[38;2;66;67;74m5[0m[38;2;79;79;86m3[0m[38;2;84;84;92mh[0m[38;2;85;85;93mh[0m[38;2;35;35;38mr[0m[38;2;2;2;2m.[0m[38;2;20;21;25m;[0m[38;2;29;30;39mr[0m[38;2;12;12;13m:[0m[38;2;21;22;29m;[0m[38;2;29;31;39mr[0m[38;2;69;69;77m5[0m[38;2;85;85;94mh[0m[38;2;84;84;92mh[0m[38;2;83;83;91mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;83;83;92mh[0m[38;2;69;69;76m5[0m[38;2;9;9;9m:[0m[38;2;182;181;180mr[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;246;246;246m#[0m[38;2;197;196;197m&[0m[38;2;232;232;232m9[0m[38;2;255;255;255mX[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m.[0m[38;2;255;255;255m;[0m[38;2;252;252;252m;[0m[38;2;251;250;250mG[0m[38;2;213;213;212mB[0m[38;2;247;246;245m9[0m[38;2;255;255;255m.[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m.[0m[38;2;255;254;251m,[0m[38;2;255;253;245mr[0m[38;2;255;252;235m2[0m[38;2;255;248;220mM[0m[38;2;255;244;205mS[0m[38;2;255;239;188mB[0m[38;2;255;230;175m&[0m[38;2;249;223;166m&[0m[38;2;255;232;180m&[0m[38;2;255;241;206mG[0m[38;2;255;247;226m5[0m[38;2;255;251;242mr[0m[38;2;255;254;253m.[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m");
    $display("[38;2;255;255;255m [0m[38;2;171;171;170m:[0m[38;2;57;60;66mX[0m[38;2;73;79;90m3[0m[38;2;198;197;197m,[0m[38;2;210;210;210m:[0m[38;2;16;15;16m;[0m[38;2;97;110;131mG[0m[38;2;154;165;187mB[0m[38;2;229;231;237m@[0m[38;2;237;240;245m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;237;239;244m@[0m[38;2;230;234;242m@[0m[38;2;89;97;111mM[0m[38;2;0;0;0m [0m[38;2;52;57;67mA[0m[38;2;128;144;171m9[0m[38;2;127;144;170m9[0m[38;2;123;138;164m#[0m[38;2;111;126;150mS[0m[38;2;113;127;151mS[0m[38;2;116;132;156m#[0m[38;2;121;137;163m#[0m[38;2;123;138;163m#[0m[38;2;27;30;36mr[0m[38;2;120;119;120mG[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;239;240;241m@[0m[38;2;203;203;208m@[0m[38;2;200;199;207m@[0m[38;2;175;172;184mB[0m[38;2;169;165;180mB[0m[38;2;170;166;180mB[0m[38;2;39;39;40mr[0m[38;2;57;57;63m2[0m[38;2;85;85;93mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;79;79;87m3[0m[38;2;67;68;75m5[0m[38;2;64;64;70m2[0m[38;2;77;77;84m3[0m[38;2;84;84;91mh[0m[38;2;84;84;92mh[0m[38;2;83;83;91mh[0m[38;2;82;82;90mh[0m[38;2;83;83;91mh[0m[38;2;70;71;78m5[0m[38;2;26;27;30mi[0m[38;2;8;8;9m,[0m[38;2;12;12;15m:[0m[38;2;10;10;13m,[0m[38;2;31;32;43mr[0m[38;2;36;37;47ms[0m[38;2;68;68;76m5[0m[38;2;84;84;91mh[0m[38;2;83;83;91mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;85;85;93mh[0m[38;2;54;54;58mA[0m[38;2;13;13;13m;[0m[38;2;203;202;201m9[0m[38;2;255;255;255mA[0m[38;2;255;255;255m [0m[38;2;255;254;254mi[0m[38;2;240;240;240m#[0m[38;2;190;190;192m&[0m[38;2;222;222;222m&[0m[38;2;255;255;255mX[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;254;254;254mi[0m[38;2;247;247;246m2[0m[38;2;252;251;251mA[0m[38;2;255;255;255m.[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m.[0m[38;2;255;255;255m.[0m[38;2;255;254;253m,[0m[38;2;255;253;250m:[0m[38;2;255;252;245mi[0m[38;2;255;250;239ms[0m[38;2;255;249;239ms[0m[38;2;255;252;246m;[0m[38;2;255;254;252m,[0m[38;2;255;255;255m:[0m[38;2;240;240;241m#[0m[38;2;220;220;220m#[0m[38;2;237;237;237mH[0m[38;2;251;251;251mX[0m[38;2;255;255;255m:[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m");
    $display("[38;2;236;236;236m#[0m[38;2;255;255;255mr[0m[38;2;220;220;219m,[0m[38;2;160;161;161mr[0m[38;2;213;213;213m;[0m[38;2;244;244;244m,[0m[38;2;50;49;49m;[0m[38;2;61;67;80m5[0m[38;2;126;143;170m9[0m[38;2;154;165;185mB[0m[38;2;230;233;238m@[0m[38;2;237;240;244m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;237;239;244m@[0m[38;2;230;234;242m@[0m[38;2;83;91;104mM[0m[38;2;0;0;0m [0m[38;2;40;43;49ms[0m[38;2;128;145;171m9[0m[38;2;100;113;133mG[0m[38;2;37;40;45ms[0m[38;2;69;69;76m5[0m[38;2;74;74;81m3[0m[38;2;66;67;74m5[0m[38;2;66;68;77m5[0m[38;2;65;69;78m5[0m[38;2;30;31;35mi[0m[38;2;72;72;73m5[0m[38;2;253;253;253m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;245;245;248m@[0m[38;2;202;200;212m@[0m[38;2;172;168;183mB[0m[38;2;132;130;141m#[0m[38;2;71;71;76m5[0m[38;2;78;78;86m3[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;78;78;85m3[0m[38;2;75;75;83m3[0m[38;2;80;80;88m3[0m[38;2;84;84;93mh[0m[38;2;83;83;92mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;84;84;92mh[0m[38;2;72;73;81m3[0m[38;2;19;20;23m;[0m[38;2;1;1;1m.[0m[38;2;28;28;29mi[0m[38;2;12;12;15m:[0m[38;2;18;19;25m;[0m[38;2;28;29;37mr[0m[38;2;52;52;59mA[0m[38;2;77;77;85m3[0m[38;2;83;83;91mh[0m[38;2;84;84;93mh[0m[38;2;84;84;93mh[0m[38;2;84;84;93mh[0m[38;2;19;20;22m;[0m[38;2;82;82;82m2[0m[38;2;188;188;189m&[0m[38;2;224;224;225m&[0m[38;2;255;255;255mi[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255ms[0m[38;2;248;248;248mA[0m[38;2;254;254;254mi[0m[38;2;251;251;250mr[0m[38;2;253;253;252mi[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255mi[0m[38;2;246;246;246m5[0m[38;2;251;251;251mA[0m[38;2;255;255;255m,[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m.[0m[38;2;248;247;247mh[0m[38;2;225;225;225m#[0m[38;2;208;208;208mB[0m[38;2;201;200;200m&[0m[38;2;206;206;207mB[0m[38;2;229;229;229m#[0m[38;2;253;253;253m2[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m");
    $display("[38;2;246;246;246mH[0m[38;2;255;255;254m;[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;248;248;248m.[0m[38;2;255;255;255m.[0m[38;2;156;156;156m;[0m[38;2;15;16;19mi[0m[38;2;113;127;151mS[0m[38;2;122;139;167m#[0m[38;2;169;178;195m&[0m[38;2;237;239;244m@[0m[38;2;236;239;244m@[0m[38;2;235;238;243m@[0m[38;2;235;238;243m@[0m[38;2;236;239;244m@[0m[38;2;232;235;243m@[0m[38;2;93;99;112mH[0m[38;2;2;2;2m.[0m[38;2;19;20;23m;[0m[38;2;113;127;150mS[0m[38;2;35;38;45ms[0m[38;2;69;68;71m5[0m[38;2;191;187;203m&[0m[38;2;188;184;200m&[0m[38;2;186;181;196m&[0m[38;2;172;169;182mB[0m[38;2;46;45;48mX[0m[38;2;3;3;2m.[0m[38;2;30;30;30mi[0m[38;2;238;238;239m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;216;216;222m@[0m[38;2;143;141;150m#[0m[38;2;89;88;94mh[0m[38;2;73;73;80m3[0m[38;2;77;77;85m3[0m[38;2;83;83;91mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;81;81;89mh[0m[38;2;83;83;91mh[0m[38;2;82;82;90mh[0m[38;2;71;71;78m5[0m[38;2;75;75;83m3[0m[38;2;85;85;93mh[0m[38;2;83;83;91mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;89mh[0m[38;2;43;44;51mX[0m[38;2;3;3;4m.[0m[38;2;70;70;74m5[0m[38;2;135;133;143m#[0m[38;2;55;54;59mA[0m[38;2;6;6;7m,[0m[38;2;8;9;10m,[0m[38;2;47;47;48mr[0m[38;2;53;53;57mX[0m[38;2;45;45;48mX[0m[38;2;49;49;53mX[0m[38;2;37;37;41mX[0m[38;2;30;30;30m;[0m[38;2;201;201;201mi[0m[38;2;255;255;255m5[0m[38;2;237;237;238m&[0m[38;2;234;233;233m&[0m[38;2;255;255;254ms[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;254;254;254mi[0m[38;2;240;239;235mG[0m[38;2;250;249;247mh[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;254;254;254mA[0m[38;2;226;226;226m&[0m[38;2;195;195;196m&[0m[38;2;215;215;215mB[0m[38;2;245;245;245mM[0m[38;2;255;255;255mi[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m:[0m[38;2;252;252;252mX[0m[38;2;240;239;239mh[0m[38;2;234;234;233mH[0m[38;2;254;254;254m2[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;252;252;252ms[0m[38;2;247;247;247mA[0m[38;2;254;254;254mr[0m[38;2;255;255;255m.[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m");
    $display("[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;251;251;251m.[0m[38;2;107;106;105m;[0m[38;2;56;62;74m5[0m[38;2;127;143;170m9[0m[38;2;123;139;166m#[0m[38;2;179;187;202m&[0m[38;2;237;240;244m@[0m[38;2;236;239;244m@[0m[38;2;235;238;243m@[0m[38;2;236;239;244m@[0m[38;2;235;238;244m@[0m[38;2;111;116;130mG[0m[38;2;14;14;15m:[0m[38;2;28;27;28m;[0m[38;2;59;64;74m2[0m[38;2;17;17;19m:[0m[38;2;128;126;134mS[0m[38;2;193;189;206m&[0m[38;2;187;183;199m&[0m[38;2;194;190;206m&[0m[38;2;114;113;120mG[0m[38;2;1;1;2m.[0m[38;2;20;21;26m;[0m[38;2;6;6;6m,[0m[38;2;136;136;137m#[0m[38;2;211;211;211m@[0m[38;2;237;237;237m@[0m[38;2;223;223;226m@[0m[38;2;135;134;141m#[0m[38;2;47;46;50mX[0m[38;2;34;34;37mr[0m[38;2;61;62;68m2[0m[38;2;74;74;81m3[0m[38;2;74;75;82m3[0m[38;2;77;77;85m3[0m[38;2;81;81;89mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;83;83;91mh[0m[38;2;35;35;39mr[0m[38;2;50;50;52mX[0m[38;2;46;46;48mX[0m[38;2;42;42;47ms[0m[38;2;78;78;85m3[0m[38;2;85;85;93mh[0m[38;2;84;84;93mh[0m[38;2;84;84;92mh[0m[38;2;84;84;93mh[0m[38;2;87;87;95mh[0m[38;2;64;65;73m5[0m[38;2;18;18;23m;[0m[38;2;13;12;12m:[0m[38;2;160;157;169mB[0m[38;2;192;188;204m&[0m[38;2;140;137;148m#[0m[38;2;63;62;66m2[0m[38;2;60;60;59mi[0m[38;2;145;144;143mH[0m[38;2;132;132;133mS[0m[38;2;192;190;186mS[0m[38;2;186;186;186m:[0m[38;2;224;224;224m,[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;251;251;251m2[0m[38;2;242;242;243mh[0m[38;2;253;252;252mr[0m[38;2;254;254;254m:[0m[38;2;254;254;254m.[0m[38;2;255;255;255m [0m[38;2;255;255;255m.[0m[38;2;255;255;255m.[0m[38;2;255;255;255m.[0m[38;2;255;255;254mr[0m[38;2;242;240;239mM[0m[38;2;252;251;251m5[0m[38;2;255;255;255m.[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m:[0m[38;2;249;249;249mh[0m[38;2;221;221;222m9[0m[38;2;196;196;197m&[0m[38;2;202;202;204m&[0m[38;2;236;236;236m#[0m[38;2;253;253;253mr[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;246;247;247mG[0m[38;2;209;208;209mB[0m[38;2;204;203;204m&[0m[38;2;214;214;214mB[0m[38;2;233;233;233mG[0m[38;2;248;247;247m5[0m");
    $display("[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;251;251;251m.[0m[38;2;134;134;135mi[0m[38;2;96;107;126mG[0m[38;2;120;137;164m9[0m[38;2;120;137;164m9[0m[38;2;171;181;198m&[0m[38;2;232;235;241m@[0m[38;2;241;243;248m@[0m[38;2;239;242;246m@[0m[38;2;242;244;249m@[0m[38;2;142;150;164m9[0m[38;2;21;22;24m:[0m[38;2;133;133;133mr[0m[38;2;28;28;29m;[0m[38;2;13;13;14m:[0m[38;2;157;154;167m9[0m[38;2;191;187;203m&[0m[38;2;188;184;200m&[0m[38;2;184;181;196m&[0m[38;2;46;46;48mX[0m[38;2;9;10;13m,[0m[38;2;33;34;44mr[0m[38;2;24;24;31mi[0m[38;2;13;14;19m:[0m[38;2;22;22;27m;[0m[38;2;37;38;41ms[0m[38;2;35;35;37mr[0m[38;2;10;10;13m,[0m[38;2;31;32;37mr[0m[38;2;57;57;64m2[0m[38;2;66;67;74m5[0m[38;2;75;75;81m3[0m[38;2;80;80;88m3[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;83;83;92mh[0m[38;2;71;71;77m5[0m[38;2;9;9;10m,[0m[38;2;178;178;179mB[0m[38;2;232;232;232m@[0m[38;2;113;112;113mG[0m[38;2;23;23;25m;[0m[38;2;49;49;53mX[0m[38;2;59;59;65m2[0m[38;2;54;54;60mA[0m[38;2;50;50;56mA[0m[38;2;52;52;56mA[0m[38;2;48;49;53mX[0m[38;2;29;30;37mr[0m[38;2;1;1;1m.[0m[38;2;100;99;104mM[0m[38;2;198;196;209m@[0m[38;2;205;202;214m@[0m[38;2;186;182;199m&[0m[38;2;141;140;149m#[0m[38;2;86;85;85mh[0m[38;2;55;55;55mA[0m[38;2;165;165;165m9[0m[38;2;255;255;255m2[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;243;243;243mS[0m[38;2;224;224;224mB[0m[38;2;255;255;254ms[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;254;254;254mA[0m[38;2;218;218;218m&[0m[38;2;187;187;187m&[0m[38;2;231;231;232m9[0m[38;2;255;255;255mX[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m.[0m[38;2;255;255;255mA[0m[38;2;232;232;232mG[0m[38;2;220;220;220m9[0m[38;2;252;252;252m5[0m[38;2;255;255;255m.[0m[38;2;255;255;255m,[0m[38;2;255;255;255m:[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m.[0m[38;2;255;255;255mi[0m[38;2;247;247;247m5[0m[38;2;232;232;232mG[0m[38;2;214;214;215mB[0m[38;2;202;202;203m&[0m");
    $display("[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;197;198;200ms[0m[38;2;157;162;171mh[0m[38;2;144;152;167mM[0m[38;2;117;129;150mG[0m[38;2;128;139;158m9[0m[38;2;167;175;189m&[0m[38;2;198;205;217m@[0m[38;2;225;229;238m@[0m[38;2;178;186;203m&[0m[38;2;35;39;47mX[0m[38;2;174;173;173m;[0m[38;2;131;131;131m;[0m[38;2;13;13;13m;[0m[38;2;167;164;176mB[0m[38;2;190;186;202m&[0m[38;2;191;187;203m&[0m[38;2;157;155;166m9[0m[38;2;12;12;12m:[0m[38;2;20;21;27m;[0m[38;2;30;31;42mr[0m[38;2;30;31;41mr[0m[38;2;31;32;42mr[0m[38;2;33;34;43mr[0m[38;2;38;39;47ms[0m[38;2;48;49;56mX[0m[38;2;67;67;75m5[0m[38;2;78;79;86m3[0m[38;2;82;82;90mh[0m[38;2;83;83;91mh[0m[38;2;83;83;91mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;85;85;93mh[0m[38;2;46;46;50mX[0m[38;2;21;21;21m;[0m[38;2;169;168;169mB[0m[38;2;203;203;203m@[0m[38;2;125;125;126mS[0m[38;2;41;40;41ms[0m[38;2;96;96;98m3[0m[38;2;24;24;24m;[0m[38;2;139;139;139m#[0m[38;2;163;163;163mB[0m[38;2;120;120;121mG[0m[38;2;6;6;5m.[0m[38;2;31;32;39mr[0m[38;2;11;12;16m:[0m[38;2;38;38;39ms[0m[38;2;181;179;191m&[0m[38;2;238;239;241m@[0m[38;2;223;222;228m@[0m[38;2;198;196;209m@[0m[38;2;236;236;239m@[0m[38;2;182;182;182m&[0m[38;2;72;72;73m3[0m[38;2;91;91;91mr[0m[38;2;212;212;213m:[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;254;253;253mi[0m[38;2;250;250;249ms[0m[38;2;249;249;249m2[0m[38;2;251;251;251mA[0m[38;2;255;255;255m.[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255mi[0m[38;2;240;240;240m#[0m[38;2;192;191;193m&[0m[38;2;200;200;201m&[0m[38;2;248;248;248mG[0m[38;2;255;255;255m:[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;254;254;254mX[0m[38;2;221;221;221m&[0m[38;2;186;186;187m9[0m[38;2;235;235;235mS[0m[38;2;255;255;255mX[0m[38;2;255;255;255m.[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m,[0m[38;2;255;255;255mr[0m");
    $display("[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m,[0m[38;2;253;253;253m2[0m[38;2;233;233;234m#[0m[38;2;203;202;203mB[0m[38;2;235;235;234mB[0m[38;2;253;253;252m;[0m[38;2;233;233;233m,[0m[38;2;188;189;191m;[0m[38;2;120;123;128mr[0m[38;2;74;78;87mA[0m[38;2;70;76;88m3[0m[38;2;94;104;122mG[0m[38;2;74;84;102mH[0m[38;2;142;142;143mi[0m[38;2;160;160;160m;[0m[38;2;24;24;24mr[0m[38;2;173;170;183mB[0m[38;2;189;185;201m&[0m[38;2;193;189;206m&[0m[38;2;126;124;134mS[0m[38;2;1;1;1m.[0m[38;2;29;30;37mr[0m[38;2;47;48;57mX[0m[38;2;56;57;65m2[0m[38;2;66;66;73m5[0m[38;2;75;75;83m3[0m[38;2;82;81;89mh[0m[38;2;84;84;92mh[0m[38;2;84;84;92mh[0m[38;2;83;83;91mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;84;84;92mh[0m[38;2;77;77;85m3[0m[38;2;72;72;79m5[0m[38;2;60;61;67m2[0m[38;2;49;49;54mX[0m[38;2;44;44;48mX[0m[38;2;18;18;20m;[0m[38;2;24;24;25m;[0m[38;2;27;27;28mi[0m[38;2;47;47;48mX[0m[38;2;181;181;182m&[0m[38;2;218;218;219m@[0m[38;2;57;56;56mA[0m[38;2;40;40;43ms[0m[38;2;54;55;62mA[0m[38;2;23;24;32mi[0m[38;2;12;12;12m:[0m[38;2;152;150;161m9[0m[38;2;228;228;233m@[0m[38;2;255;255;255m@[0m[38;2;240;239;242m@[0m[38;2;217;217;222m@[0m[38;2;255;255;255m@[0m[38;2;249;249;249m@[0m[38;2;137;137;139m#[0m[38;2;33;33;34m;[0m[38;2;213;213;213m:[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;239;239;239mB[0m[38;2;183;183;185m&[0m[38;2;246;246;246m#[0m[38;2;255;255;255m,[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m5[0m[38;2;221;221;221mB[0m[38;2;187;187;188m&[0m[38;2;221;221;221mB[0m[38;2;255;255;255m2[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;254;254;254m,[0m[38;2;250;250;249mh[0m[38;2;215;215;216m9[0m[38;2;180;180;181m&[0m[38;2;179;179;180m&[0m[38;2;220;220;221m9[0m[38;2;252;252;251m5[0m[38;2;255;255;255m,[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m");
    $display("[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255mi[0m[38;2;244;244;243mM[0m[38;2;217;217;218mB[0m[38;2;196;196;197m&[0m[38;2;208;207;208m&[0m[38;2;234;234;234mS[0m[38;2;252;252;252mA[0m[38;2;255;255;255m.[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;235;234;233m.[0m[38;2;187;186;185m,[0m[38;2;128;128;129m:[0m[38;2;94;95;97mr[0m[38;2;119;119;120ms[0m[38;2;121;121;122mr[0m[38;2;32;32;31mr[0m[38;2;183;179;192m&[0m[38;2;194;190;206m&[0m[38;2;199;195;212m@[0m[38;2;103;101;106mH[0m[38;2;0;0;0m [0m[38;2;51;51;57mA[0m[38;2;84;84;92mh[0m[38;2;84;84;92mh[0m[38;2;84;84;92mh[0m[38;2;83;83;91mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;83;83;91mh[0m[38;2;79;79;87m3[0m[38;2;39;39;43ms[0m[38;2;71;70;72m5[0m[38;2;41;41;44ms[0m[38;2;50;50;55mA[0m[38;2;81;81;89mh[0m[38;2;81;81;89mh[0m[38;2;84;84;92mh[0m[38;2;75;75;83m3[0m[38;2;70;70;77m5[0m[38;2;54;54;60mA[0m[38;2;24;24;26mi[0m[38;2;24;24;26mi[0m[38;2;38;38;42ms[0m[38;2;85;85;93mh[0m[38;2;64;64;72m2[0m[38;2;27;28;37mi[0m[38;2;5;5;5m.[0m[38;2;120;120;130mS[0m[38;2;216;214;224m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;248;249;249m@[0m[38;2;240;241;243m@[0m[38;2;255;255;255m@[0m[38;2;186;186;188m&[0m[38;2;19;18;18m;[0m[38;2;210;210;210m:[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255ms[0m[38;2;225;225;226mB[0m[38;2;176;176;177m&[0m[38;2;241;241;241m9[0m[38;2;255;255;255m;[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m:[0m[38;2;247;247;247mH[0m[38;2;202;201;202m&[0m[38;2;192;192;193m&[0m[38;2;241;241;241mS[0m[38;2;255;255;255mi[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m.[0m[38;2;255;255;255mA[0m[38;2;231;232;232mS[0m[38;2;198;198;198mB[0m[38;2;193;193;194m&[0m[38;2;216;216;216mB[0m[38;2;246;246;246mM[0m[38;2;255;255;255mi[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m");
    $display("[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;248;248;248mG[0m[38;2;205;205;206m&[0m[38;2;198;197;198m&[0m[38;2;221;221;222m9[0m[38;2;248;248;248m3[0m[38;2;255;255;255m;[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m.[0m[38;2;221;221;221m,[0m[38;2;112;113;112m;[0m[38;2;22;22;22mi[0m[38;2;137;134;144m#[0m[38;2;137;134;146m#[0m[38;2;130;128;138mS[0m[38;2;64;63;65m2[0m[38;2;5;6;7m,[0m[38;2;71;72;79m5[0m[38;2;83;83;92mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;83;83;91mh[0m[38;2;73;74;80m3[0m[38;2;5;5;5m.[0m[38;2;169;169;170mB[0m[38;2;221;221;222m@[0m[38;2;89;89;90mh[0m[38;2;21;21;22m;[0m[38;2;57;56;59mA[0m[38;2;27;27;30mi[0m[38;2;43;43;46ms[0m[38;2;66;66;68m2[0m[38;2;77;77;79m3[0m[38;2;16;16;16m:[0m[38;2;43;44;48mX[0m[38;2;87;87;96mh[0m[38;2;82;82;90mh[0m[38;2;57;57;65m2[0m[38;2;27;28;35mi[0m[38;2;4;4;4m.[0m[38;2;127;126;136mS[0m[38;2;208;206;216m@[0m[38;2;255;255;254m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;243;243;243m@[0m[38;2;55;55;56m2[0m[38;2;110;109;109m:[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255mi[0m[38;2;232;232;232mB[0m[38;2;174;174;175m&[0m[38;2;235;235;235m9[0m[38;2;255;255;255mi[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255mX[0m[38;2;231;231;232m9[0m[38;2;187;187;188m&[0m[38;2;230;230;230m&[0m[38;2;255;255;255mi[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m;[0m[38;2;248;248;248m3[0m[38;2;221;221;222m9[0m[38;2;198;198;199m&[0m[38;2;204;204;205m&[0m[38;2;236;236;236mS[0m[38;2;254;254;254mX[0m[38;2;254;254;254m.[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m");
    $display("[38;2;242;242;241mH[0m[38;2;236;236;236mG[0m[38;2;254;254;254mi[0m[38;2;251;251;251mA[0m[38;2;240;240;241m5[0m[38;2;255;255;255ms[0m[38;2;255;255;255m.[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m.[0m[38;2;125;126;125m;[0m[38;2;54;54;55ms[0m[38;2;91;89;96mh[0m[38;2;88;86;93mh[0m[38;2;98;96;103mM[0m[38;2;105;103;110mH[0m[38;2;118;116;125mG[0m[38;2;96;95;102mM[0m[38;2;7;7;8m,[0m[38;2;73;73;80m3[0m[38;2;84;83;92mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;84;84;93mh[0m[38;2;59;60;65m2[0m[38;2;12;11;12m,[0m[38;2;184;184;185m&[0m[38;2;211;211;211m@[0m[38;2;115;115;115mG[0m[38;2;30;29;29mi[0m[38;2;129;129;131mS[0m[38;2;39;38;39ms[0m[38;2;204;204;204m@[0m[38;2;253;253;253m@[0m[38;2;142;141;143m#[0m[38;2;15;15;16m:[0m[38;2;71;71;77m5[0m[38;2;67;67;75m5[0m[38;2;42;43;51mX[0m[38;2;30;31;41mr[0m[38;2;13;13;16m:[0m[38;2;47;47;49mX[0m[38;2;176;172;187m&[0m[38;2;200;198;209m@[0m[38;2;254;255;254m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;106;106;106mG[0m[38;2;56;56;56m:[0m[38;2;237;237;237mM[0m[38;2;232;232;233mG[0m[38;2;255;255;255mA[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m;[0m[38;2;239;239;239m9[0m[38;2;178;177;179m&[0m[38;2;240;240;240mB[0m[38;2;255;255;255m.[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m.[0m[38;2;251;251;251mA[0m[38;2;246;246;246m2[0m[38;2;254;254;254m,[0m[38;2;255;255;255m.[0m[38;2;255;255;255m.[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m.[0m[38;2;255;255;255mA[0m[38;2;234;234;234mS[0m[38;2;202;202;203m&[0m[38;2;218;218;219m&[0m[38;2;254;254;254m5[0m[38;2;255;255;255m,[0m[38;2;255;255;255m:[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m");
    $display("[38;2;229;229;229m#[0m[38;2;233;233;233m#[0m[38;2;254;254;254mi[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m,[0m[38;2;93;93;93ms[0m[38;2;55;54;56m2[0m[38;2;234;233;239m@[0m[38;2;240;239;244m@[0m[38;2;243;242;247m@[0m[38;2;246;245;249m@[0m[38;2;248;248;251m@[0m[38;2;216;216;221m@[0m[38;2;35;35;37mr[0m[38;2;32;32;35mr[0m[38;2;85;85;93mh[0m[38;2;83;83;91mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;83;83;91mh[0m[38;2;69;69;76m5[0m[38;2;35;35;38mr[0m[38;2;48;48;50mX[0m[38;2;45;45;49mX[0m[38;2;48;48;52mX[0m[38;2;51;51;55mA[0m[38;2;47;47;52mX[0m[38;2;52;51;53mA[0m[38;2;106;106;107mH[0m[38;2;126;126;128mS[0m[38;2;19;18;19m;[0m[38;2;44;44;49mX[0m[38;2;45;46;55mX[0m[38;2;31;32;42mr[0m[38;2;27;28;37mi[0m[38;2;12;13;16m:[0m[38;2;29;29;30mi[0m[38;2;162;159;171mB[0m[38;2;191;187;204m&[0m[38;2;189;185;200m&[0m[38;2;239;238;240m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;134;134;135m#[0m[38;2;37;37;38m:[0m[38;2;216;216;217m,[0m[38;2;255;255;255mH[0m[38;2;173;172;174m&[0m[38;2;232;232;233mB[0m[38;2;255;255;255m:[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m:[0m[38;2;247;247;248m3[0m[38;2;240;240;240mB[0m[38;2;231;230;231mS[0m[38;2;255;255;255mX[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m.[0m[38;2;245;245;245m#[0m[38;2;218;217;217mB[0m[38;2;254;254;254m3[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m;[0m[38;2;253;253;253mi[0m[38;2;254;254;254m2[0m[38;2;217;217;218m&[0m[38;2;189;189;190m9[0m[38;2;236;235;236mS[0m[38;2;255;255;255mX[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m");
    $display("[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m,[0m[38;2;243;243;243mB[0m[38;2;149;148;148m9[0m[38;2;19;19;19m;[0m[38;2;193;193;194m&[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;182;182;185m&[0m[38;2;31;31;31mi[0m[38;2;34;34;37mr[0m[38;2;79;80;87m3[0m[38;2;85;85;93mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;83;83;91mh[0m[38;2;84;84;92mh[0m[38;2;82;82;90mh[0m[38;2;83;83;92mh[0m[38;2;85;85;93mh[0m[38;2;85;85;93mh[0m[38;2;85;85;93mh[0m[38;2;81;81;88mh[0m[38;2;57;57;63m2[0m[38;2;24;24;30mi[0m[38;2;27;27;35mi[0m[38;2;34;34;45ms[0m[38;2;26;27;36mi[0m[38;2;12;13;17m:[0m[38;2;16;16;17m:[0m[38;2;92;92;99mM[0m[38;2;47;47;50mX[0m[38;2;104;102;109mH[0m[38;2;194;190;206m&[0m[38;2;186;181;198m&[0m[38;2;201;200;210m@[0m[38;2;250;250;252m@[0m[38;2;135;134;135m#[0m[38;2;39;38;38m;[0m[38;2;204;204;204m:[0m[38;2;255;255;255m [0m[38;2;255;255;255m:[0m[38;2;233;233;234mB[0m[38;2;172;172;173m&[0m[38;2;254;254;254mG[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;249;249;249mS[0m[38;2;185;185;186m&[0m[38;2;213;213;214m&[0m[38;2;255;255;255m2[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;251;251;251m2[0m[38;2;239;239;239mM[0m[38;2;255;254;255mX[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m,[0m[38;2;248;248;248mh[0m[38;2;216;216;216m9[0m[38;2;178;178;178m&[0m[38;2;181;181;182m&[0m[38;2;222;222;222m9[0m[38;2;251;250;250m3[0m[38;2;254;254;254m,[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m");
    $display("[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;254;254;254m:[0m[38;2;252;252;252mr[0m[38;2;253;253;253mr[0m[38;2;242;242;242mM[0m[38;2;239;239;239mh[0m[38;2;109;109;108mr[0m[38;2;57;57;58m5[0m[38;2;243;244;244m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;219;219;219m@[0m[38;2;87;87;89mh[0m[38;2;28;28;29mi[0m[38;2;53;53;59mA[0m[38;2;81;81;90mh[0m[38;2;85;85;93mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;83;83;91mh[0m[38;2;84;84;92mh[0m[38;2;77;77;85m3[0m[38;2;60;60;68m2[0m[38;2;41;42;52mX[0m[38;2;30;31;41mr[0m[38;2;20;21;28m;[0m[38;2;9;9;13m,[0m[38;2;13;12;14m:[0m[38;2;58;57;61mA[0m[38;2;150;149;157m9[0m[38;2;233;233;239m@[0m[38;2;183;182;184m&[0m[38;2;27;26;26mi[0m[38;2;131;129;138mS[0m[38;2;197;193;210m&[0m[38;2;177;174;189m&[0m[38;2;89;89;93mM[0m[38;2;58;58;57m;[0m[38;2;211;211;210m:[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m3[0m[38;2;188;188;189m&[0m[38;2;208;208;209m&[0m[38;2;255;255;255ms[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m.[0m[38;2;252;252;252mG[0m[38;2;187;186;187m&[0m[38;2;206;206;207m&[0m[38;2;255;255;255m3[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;254;254;254mr[0m[38;2;250;250;251mA[0m[38;2;255;255;255mi[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m.[0m[38;2;255;255;255mA[0m[38;2;233;233;233mS[0m[38;2;189;189;189mB[0m[38;2;209;209;210m&[0m[38;2;253;253;252m3[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m");
    $display("[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m,[0m[38;2;242;242;242m9[0m[38;2;203;202;203m&[0m[38;2;253;253;252mG[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;242;242;242m,[0m[38;2;96;96;96m:[0m[38;2;69;69;70m5[0m[38;2;179;179;180m&[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;200;200;201m&[0m[38;2;111;110;113mH[0m[38;2;34;33;36mr[0m[38;2;53;53;58mA[0m[38;2;81;81;89mh[0m[38;2;85;85;93mh[0m[38;2;83;83;91mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;82;82;90mh[0m[38;2;83;83;91mh[0m[38;2;84;84;92mh[0m[38;2;83;83;91mh[0m[38;2;73;74;81m3[0m[38;2;51;52;60mA[0m[38;2;28;29;37mr[0m[38;2;15;16;22m:[0m[38;2;13;14;18m:[0m[38;2;24;25;28mi[0m[38;2;54;54;58mA[0m[38;2;102;101;109mH[0m[38;2;168;167;175mB[0m[38;2;229;228;234m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;169;169;170mB[0m[38;2;28;27;28mi[0m[38;2;122;119;128mS[0m[38;2;101;100;105m5[0m[38;2;129;129;129m:[0m[38;2;238;238;238m,[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m.[0m[38;2;247;247;247m9[0m[38;2;166;165;167mB[0m[38;2;247;247;247m9[0m[38;2;255;255;255m.[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;254;254;254mM[0m[38;2;194;193;195m&[0m[38;2;197;197;198m&[0m[38;2;255;255;255mh[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;252;252;252mG[0m[38;2;198;197;199m&[0m[38;2;226;226;226m&[0m[38;2;254;254;254ms[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m:[0m[38;2;253;253;253m;[0m[38;2;254;254;254m,[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m");
    $display("[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m.[0m[38;2;253;252;252ms[0m[38;2;252;251;250mX[0m[38;2;255;255;254m:[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m.[0m[38;2;188;187;188m,[0m[38;2;57;57;58m;[0m[38;2;106;105;107mG[0m[38;2;236;236;237m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;186;185;186m&[0m[38;2;70;70;71m5[0m[38;2;30;30;32mi[0m[38;2;47;47;52mX[0m[38;2;69;69;76m5[0m[38;2;80;80;87m3[0m[38;2;83;83;92mh[0m[38;2;84;84;93mh[0m[38;2;84;85;93mh[0m[38;2;84;84;93mh[0m[38;2;84;84;93mh[0m[38;2;84;84;92mh[0m[38;2;82;82;90mh[0m[38;2;75;76;83m3[0m[38;2;59;59;65m2[0m[38;2;37;38;43ms[0m[38;2;20;21;25m;[0m[38;2;18;18;22m;[0m[38;2;47;47;52mX[0m[38;2;88;87;94mh[0m[38;2;132;129;139mS[0m[38;2;167;164;178mB[0m[38;2;201;198;210m@[0m[38;2;234;233;239m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;151;151;153m9[0m[38;2;13;13;14m,[0m[38;2;204;204;203m:[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255mr[0m[38;2;213;213;213m&[0m[38;2;188;188;189m&[0m[38;2;255;255;255m3[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255mh[0m[38;2;202;202;203m&[0m[38;2;192;192;193m&[0m[38;2;254;253;253mH[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m,[0m[38;2;249;249;249mA[0m[38;2;243;243;243m2[0m[38;2;254;254;254m;[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m");
    $display("[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m:[0m[38;2;249;249;249mH[0m[38;2;213;213;213mS[0m[38;2;248;248;248mH[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;237;237;237m,[0m[38;2;113;113;113m:[0m[38;2;62;62;63m2[0m[38;2;169;169;170mB[0m[38;2;244;244;244m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;253;254;254m@[0m[38;2;191;191;194m&[0m[38;2;108;107;113mH[0m[38;2;62;61;65m2[0m[38;2;47;47;50mX[0m[38;2;46;46;50mX[0m[38;2;48;48;52mX[0m[38;2;50;50;54mX[0m[38;2;51;51;55mA[0m[38;2;49;49;53mX[0m[38;2;45;45;49mX[0m[38;2;38;38;42ms[0m[38;2;41;41;44ms[0m[38;2;57;57;60mA[0m[38;2;44;44;45ms[0m[38;2;25;25;26mi[0m[38;2;129;127;136mS[0m[38;2;190;186;202m&[0m[38;2;197;193;210m&[0m[38;2;205;202;216m@[0m[38;2;236;235;241m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;255;255;255m@[0m[38;2;245;245;245m@[0m[38;2;232;232;232m@[0m[38;2;208;208;209m@[0m[38;2;162;162;163mB[0m[38;2;97;97;98mM[0m[38;2;49;48;49mA[0m[38;2;223;222;221mG[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255mH[0m[38;2;176;175;176m&[0m[38;2;229;228;228mB[0m[38;2;255;255;255m:[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m5[0m[38;2;210;210;211m&[0m[38;2;189;188;189m&[0m[38;2;250;250;250mS[0m[38;2;255;255;255m,[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;254;254;254m.[0m[38;2;255;255;255m:[0m[38;2;255;255;255m.[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m");
    $display("[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;254;254;254ms[0m[38;2;233;233;234mB[0m[38;2;184;183;184m&[0m[38;2;213;213;213m&[0m[38;2;252;252;252m3[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m.[0m[38;2;191;191;191m,[0m[38;2;89;89;89m;[0m[38;2;75;75;76m5[0m[38;2;133;133;134m#[0m[38;2;188;188;189m&[0m[38;2;220;220;221m@[0m[38;2;234;233;234m@[0m[38;2;240;240;241m@[0m[38;2;244;244;245m@[0m[38;2;246;246;246m@[0m[38;2;231;231;233m@[0m[38;2;182;180;190m&[0m[38;2;149;147;158m9[0m[38;2;135;132;142m#[0m[38;2;130;128;137mS[0m[38;2;123;121;130mS[0m[38;2;122;120;129mS[0m[38;2;128;126;135mS[0m[38;2;142;139;151m#[0m[38;2;143;141;153m#[0m[38;2;115;114;122mG[0m[38;2;75;74;78m3[0m[38;2;41;41;41mr[0m[38;2;47;46;46mX[0m[38;2;68;68;70m5[0m[38;2;79;78;83m3[0m[38;2;94;93;100mM[0m[38;2;133;133;136m#[0m[38;2;161;161;161mB[0m[38;2;154;154;156m9[0m[38;2;141;141;141m#[0m[38;2;122;122;123mS[0m[38;2;97;97;97mM[0m[38;2;92;91;92m5[0m[38;2;113;113;113ms[0m[38;2;111;111;111mi[0m[38;2;135;135;136m,[0m[38;2;199;199;199m2[0m[38;2;172;171;172mB[0m[38;2;229;229;229mB[0m[38;2;255;255;255m,[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m:[0m[38;2;241;241;241mS[0m[38;2;234;234;234mS[0m[38;2;255;255;255m;[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m2[0m[38;2;213;213;214m&[0m[38;2;182;182;183m&[0m[38;2;250;250;250mS[0m[38;2;255;255;255m.[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;254;254;254mX[0m[38;2;218;218;219mB[0m[38;2;230;230;230m9[0m[38;2;254;254;254mX[0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m[38;2;255;255;255m [0m");
	$display("\033[0;32m \033[5m    //   ) )     // | |     //   ) )     //   ) )\033[m");
    $display("\033[0;32m \033[5m   //___/ /     //__| |    ((           ((\033[m");
    $display("\033[0;32m \033[5m  / ____ /     / ___  |      \\           \\\033[m");
    $display("\033[0;32m \033[5m //           //    | |        ) )          ) )\033[m");
    $display("\033[0;32m \033[5m//           //     | | ((___ / /    ((___ / /\033[m");
	$display("**************************************************");
	$display("                  Congratulations!                ");
	$display("              execution cycles = %7d", total_latency);
	$display("              clock period = %4fns", CYCLE);
	$display("**************************************************");
end endtask
endmodule
